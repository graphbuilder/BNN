module test_layer_all(
clk, 
rstn
);
input clk;
input rstn;

wire P0000;
wire P0010;
wire P0020;
wire P0030;
wire P0040;
wire P0050;
wire P0060;
wire P0070;
wire P0080;
wire P0090;
wire P00A0;
wire P00B0;
wire P00C0;
wire P00D0;
wire P00E0;
wire P00F0;
wire P0100;
wire P0110;
wire P0120;
wire P0130;
wire P0140;
wire P0150;
wire P0160;
wire P0170;
wire P0180;
wire P0190;
wire P01A0;
wire P01B0;
wire P01C0;
wire P01D0;
wire P01E0;
wire P01F0;
wire P0200;
wire P0210;
wire P0220;
wire P0230;
wire P0240;
wire P0250;
wire P0260;
wire P0270;
wire P0280;
wire P0290;
wire P02A0;
wire P02B0;
wire P02C0;
wire P02D0;
wire P02E0;
wire P02F0;
wire P0300;
wire P0310;
wire P0320;
wire P0330;
wire P0340;
wire P0350;
wire P0360;
wire P0370;
wire P0380;
wire P0390;
wire P03A0;
wire P03B0;
wire P03C0;
wire P03D0;
wire P03E0;
wire P03F0;
wire P0400;
wire P0410;
wire P0420;
wire P0430;
wire P0440;
wire P0450;
wire P0460;
wire P0470;
wire P0480;
wire P0490;
wire P04A0;
wire P04B0;
wire P04C0;
wire P04D0;
wire P04E0;
wire P04F0;
wire P0500;
wire P0510;
wire P0520;
wire P0530;
wire P0540;
wire P0550;
wire P0560;
wire P0570;
wire P0580;
wire P0590;
wire P05A0;
wire P05B0;
wire P05C0;
wire P05D0;
wire P05E0;
wire P05F0;
wire P0600;
wire P0610;
wire P0620;
wire P0630;
wire P0640;
wire P0650;
wire P0660;
wire P0670;
wire P0680;
wire P0690;
wire P06A0;
wire P06B0;
wire P06C0;
wire P06D0;
wire P06E0;
wire P06F0;
wire P0700;
wire P0710;
wire P0720;
wire P0730;
wire P0740;
wire P0750;
wire P0760;
wire P0770;
wire P0780;
wire P0790;
wire P07A0;
wire P07B0;
wire P07C0;
wire P07D0;
wire P07E0;
wire P07F0;
wire P0800;
wire P0810;
wire P0820;
wire P0830;
wire P0840;
wire P0850;
wire P0860;
wire P0870;
wire P0880;
wire P0890;
wire P08A0;
wire P08B0;
wire P08C0;
wire P08D0;
wire P08E0;
wire P08F0;
wire P0900;
wire P0910;
wire P0920;
wire P0930;
wire P0940;
wire P0950;
wire P0960;
wire P0970;
wire P0980;
wire P0990;
wire P09A0;
wire P09B0;
wire P09C0;
wire P09D0;
wire P09E0;
wire P09F0;
wire P0A00;
wire P0A10;
wire P0A20;
wire P0A30;
wire P0A40;
wire P0A50;
wire P0A60;
wire P0A70;
wire P0A80;
wire P0A90;
wire P0AA0;
wire P0AB0;
wire P0AC0;
wire P0AD0;
wire P0AE0;
wire P0AF0;
wire P0B00;
wire P0B10;
wire P0B20;
wire P0B30;
wire P0B40;
wire P0B50;
wire P0B60;
wire P0B70;
wire P0B80;
wire P0B90;
wire P0BA0;
wire P0BB0;
wire P0BC0;
wire P0BD0;
wire P0BE0;
wire P0BF0;
wire P0C00;
wire P0C10;
wire P0C20;
wire P0C30;
wire P0C40;
wire P0C50;
wire P0C60;
wire P0C70;
wire P0C80;
wire P0C90;
wire P0CA0;
wire P0CB0;
wire P0CC0;
wire P0CD0;
wire P0CE0;
wire P0CF0;
wire P0D00;
wire P0D10;
wire P0D20;
wire P0D30;
wire P0D40;
wire P0D50;
wire P0D60;
wire P0D70;
wire P0D80;
wire P0D90;
wire P0DA0;
wire P0DB0;
wire P0DC0;
wire P0DD0;
wire P0DE0;
wire P0DF0;
wire P0E00;
wire P0E10;
wire P0E20;
wire P0E30;
wire P0E40;
wire P0E50;
wire P0E60;
wire P0E70;
wire P0E80;
wire P0E90;
wire P0EA0;
wire P0EB0;
wire P0EC0;
wire P0ED0;
wire P0EE0;
wire P0EF0;
wire P0F00;
wire P0F10;
wire P0F20;
wire P0F30;
wire P0F40;
wire P0F50;
wire P0F60;
wire P0F70;
wire P0F80;
wire P0F90;
wire P0FA0;
wire P0FB0;
wire P0FC0;
wire P0FD0;
wire P0FE0;
wire P0FF0;
wire P0001;
wire P0011;
wire P0021;
wire P0031;
wire P0041;
wire P0051;
wire P0061;
wire P0071;
wire P0081;
wire P0091;
wire P00A1;
wire P00B1;
wire P00C1;
wire P00D1;
wire P00E1;
wire P00F1;
wire P0101;
wire P0111;
wire P0121;
wire P0131;
wire P0141;
wire P0151;
wire P0161;
wire P0171;
wire P0181;
wire P0191;
wire P01A1;
wire P01B1;
wire P01C1;
wire P01D1;
wire P01E1;
wire P01F1;
wire P0201;
wire P0211;
wire P0221;
wire P0231;
wire P0241;
wire P0251;
wire P0261;
wire P0271;
wire P0281;
wire P0291;
wire P02A1;
wire P02B1;
wire P02C1;
wire P02D1;
wire P02E1;
wire P02F1;
wire P0301;
wire P0311;
wire P0321;
wire P0331;
wire P0341;
wire P0351;
wire P0361;
wire P0371;
wire P0381;
wire P0391;
wire P03A1;
wire P03B1;
wire P03C1;
wire P03D1;
wire P03E1;
wire P03F1;
wire P0401;
wire P0411;
wire P0421;
wire P0431;
wire P0441;
wire P0451;
wire P0461;
wire P0471;
wire P0481;
wire P0491;
wire P04A1;
wire P04B1;
wire P04C1;
wire P04D1;
wire P04E1;
wire P04F1;
wire P0501;
wire P0511;
wire P0521;
wire P0531;
wire P0541;
wire P0551;
wire P0561;
wire P0571;
wire P0581;
wire P0591;
wire P05A1;
wire P05B1;
wire P05C1;
wire P05D1;
wire P05E1;
wire P05F1;
wire P0601;
wire P0611;
wire P0621;
wire P0631;
wire P0641;
wire P0651;
wire P0661;
wire P0671;
wire P0681;
wire P0691;
wire P06A1;
wire P06B1;
wire P06C1;
wire P06D1;
wire P06E1;
wire P06F1;
wire P0701;
wire P0711;
wire P0721;
wire P0731;
wire P0741;
wire P0751;
wire P0761;
wire P0771;
wire P0781;
wire P0791;
wire P07A1;
wire P07B1;
wire P07C1;
wire P07D1;
wire P07E1;
wire P07F1;
wire P0801;
wire P0811;
wire P0821;
wire P0831;
wire P0841;
wire P0851;
wire P0861;
wire P0871;
wire P0881;
wire P0891;
wire P08A1;
wire P08B1;
wire P08C1;
wire P08D1;
wire P08E1;
wire P08F1;
wire P0901;
wire P0911;
wire P0921;
wire P0931;
wire P0941;
wire P0951;
wire P0961;
wire P0971;
wire P0981;
wire P0991;
wire P09A1;
wire P09B1;
wire P09C1;
wire P09D1;
wire P09E1;
wire P09F1;
wire P0A01;
wire P0A11;
wire P0A21;
wire P0A31;
wire P0A41;
wire P0A51;
wire P0A61;
wire P0A71;
wire P0A81;
wire P0A91;
wire P0AA1;
wire P0AB1;
wire P0AC1;
wire P0AD1;
wire P0AE1;
wire P0AF1;
wire P0B01;
wire P0B11;
wire P0B21;
wire P0B31;
wire P0B41;
wire P0B51;
wire P0B61;
wire P0B71;
wire P0B81;
wire P0B91;
wire P0BA1;
wire P0BB1;
wire P0BC1;
wire P0BD1;
wire P0BE1;
wire P0BF1;
wire P0C01;
wire P0C11;
wire P0C21;
wire P0C31;
wire P0C41;
wire P0C51;
wire P0C61;
wire P0C71;
wire P0C81;
wire P0C91;
wire P0CA1;
wire P0CB1;
wire P0CC1;
wire P0CD1;
wire P0CE1;
wire P0CF1;
wire P0D01;
wire P0D11;
wire P0D21;
wire P0D31;
wire P0D41;
wire P0D51;
wire P0D61;
wire P0D71;
wire P0D81;
wire P0D91;
wire P0DA1;
wire P0DB1;
wire P0DC1;
wire P0DD1;
wire P0DE1;
wire P0DF1;
wire P0E01;
wire P0E11;
wire P0E21;
wire P0E31;
wire P0E41;
wire P0E51;
wire P0E61;
wire P0E71;
wire P0E81;
wire P0E91;
wire P0EA1;
wire P0EB1;
wire P0EC1;
wire P0ED1;
wire P0EE1;
wire P0EF1;
wire P0F01;
wire P0F11;
wire P0F21;
wire P0F31;
wire P0F41;
wire P0F51;
wire P0F61;
wire P0F71;
wire P0F81;
wire P0F91;
wire P0FA1;
wire P0FB1;
wire P0FC1;
wire P0FD1;
wire P0FE1;
wire P0FF1;
wire P0002;
wire P0012;
wire P0022;
wire P0032;
wire P0042;
wire P0052;
wire P0062;
wire P0072;
wire P0082;
wire P0092;
wire P00A2;
wire P00B2;
wire P00C2;
wire P00D2;
wire P00E2;
wire P00F2;
wire P0102;
wire P0112;
wire P0122;
wire P0132;
wire P0142;
wire P0152;
wire P0162;
wire P0172;
wire P0182;
wire P0192;
wire P01A2;
wire P01B2;
wire P01C2;
wire P01D2;
wire P01E2;
wire P01F2;
wire P0202;
wire P0212;
wire P0222;
wire P0232;
wire P0242;
wire P0252;
wire P0262;
wire P0272;
wire P0282;
wire P0292;
wire P02A2;
wire P02B2;
wire P02C2;
wire P02D2;
wire P02E2;
wire P02F2;
wire P0302;
wire P0312;
wire P0322;
wire P0332;
wire P0342;
wire P0352;
wire P0362;
wire P0372;
wire P0382;
wire P0392;
wire P03A2;
wire P03B2;
wire P03C2;
wire P03D2;
wire P03E2;
wire P03F2;
wire P0402;
wire P0412;
wire P0422;
wire P0432;
wire P0442;
wire P0452;
wire P0462;
wire P0472;
wire P0482;
wire P0492;
wire P04A2;
wire P04B2;
wire P04C2;
wire P04D2;
wire P04E2;
wire P04F2;
wire P0502;
wire P0512;
wire P0522;
wire P0532;
wire P0542;
wire P0552;
wire P0562;
wire P0572;
wire P0582;
wire P0592;
wire P05A2;
wire P05B2;
wire P05C2;
wire P05D2;
wire P05E2;
wire P05F2;
wire P0602;
wire P0612;
wire P0622;
wire P0632;
wire P0642;
wire P0652;
wire P0662;
wire P0672;
wire P0682;
wire P0692;
wire P06A2;
wire P06B2;
wire P06C2;
wire P06D2;
wire P06E2;
wire P06F2;
wire P0702;
wire P0712;
wire P0722;
wire P0732;
wire P0742;
wire P0752;
wire P0762;
wire P0772;
wire P0782;
wire P0792;
wire P07A2;
wire P07B2;
wire P07C2;
wire P07D2;
wire P07E2;
wire P07F2;
wire P0802;
wire P0812;
wire P0822;
wire P0832;
wire P0842;
wire P0852;
wire P0862;
wire P0872;
wire P0882;
wire P0892;
wire P08A2;
wire P08B2;
wire P08C2;
wire P08D2;
wire P08E2;
wire P08F2;
wire P0902;
wire P0912;
wire P0922;
wire P0932;
wire P0942;
wire P0952;
wire P0962;
wire P0972;
wire P0982;
wire P0992;
wire P09A2;
wire P09B2;
wire P09C2;
wire P09D2;
wire P09E2;
wire P09F2;
wire P0A02;
wire P0A12;
wire P0A22;
wire P0A32;
wire P0A42;
wire P0A52;
wire P0A62;
wire P0A72;
wire P0A82;
wire P0A92;
wire P0AA2;
wire P0AB2;
wire P0AC2;
wire P0AD2;
wire P0AE2;
wire P0AF2;
wire P0B02;
wire P0B12;
wire P0B22;
wire P0B32;
wire P0B42;
wire P0B52;
wire P0B62;
wire P0B72;
wire P0B82;
wire P0B92;
wire P0BA2;
wire P0BB2;
wire P0BC2;
wire P0BD2;
wire P0BE2;
wire P0BF2;
wire P0C02;
wire P0C12;
wire P0C22;
wire P0C32;
wire P0C42;
wire P0C52;
wire P0C62;
wire P0C72;
wire P0C82;
wire P0C92;
wire P0CA2;
wire P0CB2;
wire P0CC2;
wire P0CD2;
wire P0CE2;
wire P0CF2;
wire P0D02;
wire P0D12;
wire P0D22;
wire P0D32;
wire P0D42;
wire P0D52;
wire P0D62;
wire P0D72;
wire P0D82;
wire P0D92;
wire P0DA2;
wire P0DB2;
wire P0DC2;
wire P0DD2;
wire P0DE2;
wire P0DF2;
wire P0E02;
wire P0E12;
wire P0E22;
wire P0E32;
wire P0E42;
wire P0E52;
wire P0E62;
wire P0E72;
wire P0E82;
wire P0E92;
wire P0EA2;
wire P0EB2;
wire P0EC2;
wire P0ED2;
wire P0EE2;
wire P0EF2;
wire P0F02;
wire P0F12;
wire P0F22;
wire P0F32;
wire P0F42;
wire P0F52;
wire P0F62;
wire P0F72;
wire P0F82;
wire P0F92;
wire P0FA2;
wire P0FB2;
wire P0FC2;
wire P0FD2;
wire P0FE2;
wire P0FF2;
wire P1000;
wire P1010;
wire P1020;
wire P1030;
wire P1040;
wire P1050;
wire P1060;
wire P1100;
wire P1110;
wire P1120;
wire P1130;
wire P1140;
wire P1150;
wire P1160;
wire P1200;
wire P1210;
wire P1220;
wire P1230;
wire P1240;
wire P1250;
wire P1260;
wire P1300;
wire P1310;
wire P1320;
wire P1330;
wire P1340;
wire P1350;
wire P1360;
wire P1400;
wire P1410;
wire P1420;
wire P1430;
wire P1440;
wire P1450;
wire P1460;
wire P1500;
wire P1510;
wire P1520;
wire P1530;
wire P1540;
wire P1550;
wire P1560;
wire P1600;
wire P1610;
wire P1620;
wire P1630;
wire P1640;
wire P1650;
wire P1660;
wire P1001;
wire P1011;
wire P1021;
wire P1031;
wire P1041;
wire P1051;
wire P1061;
wire P1101;
wire P1111;
wire P1121;
wire P1131;
wire P1141;
wire P1151;
wire P1161;
wire P1201;
wire P1211;
wire P1221;
wire P1231;
wire P1241;
wire P1251;
wire P1261;
wire P1301;
wire P1311;
wire P1321;
wire P1331;
wire P1341;
wire P1351;
wire P1361;
wire P1401;
wire P1411;
wire P1421;
wire P1431;
wire P1441;
wire P1451;
wire P1461;
wire P1501;
wire P1511;
wire P1521;
wire P1531;
wire P1541;
wire P1551;
wire P1561;
wire P1601;
wire P1611;
wire P1621;
wire P1631;
wire P1641;
wire P1651;
wire P1661;
wire P1002;
wire P1012;
wire P1022;
wire P1032;
wire P1042;
wire P1052;
wire P1062;
wire P1102;
wire P1112;
wire P1122;
wire P1132;
wire P1142;
wire P1152;
wire P1162;
wire P1202;
wire P1212;
wire P1222;
wire P1232;
wire P1242;
wire P1252;
wire P1262;
wire P1302;
wire P1312;
wire P1322;
wire P1332;
wire P1342;
wire P1352;
wire P1362;
wire P1402;
wire P1412;
wire P1422;
wire P1432;
wire P1442;
wire P1452;
wire P1462;
wire P1502;
wire P1512;
wire P1522;
wire P1532;
wire P1542;
wire P1552;
wire P1562;
wire P1602;
wire P1612;
wire P1622;
wire P1632;
wire P1642;
wire P1652;
wire P1662;
wire W00000,W00010,W00020,W00100,W00110,W00120,W00200,W00210,W00220;
wire W00001,W00011,W00021,W00101,W00111,W00121,W00201,W00211,W00221;
wire W00002,W00012,W00022,W00102,W00112,W00122,W00202,W00212,W00222;
wire W01000,W01010,W01020,W01100,W01110,W01120,W01200,W01210,W01220;
wire W01001,W01011,W01021,W01101,W01111,W01121,W01201,W01211,W01221;
wire W01002,W01012,W01022,W01102,W01112,W01122,W01202,W01212,W01222;
wire W02000,W02010,W02020,W02100,W02110,W02120,W02200,W02210,W02220;
wire W02001,W02011,W02021,W02101,W02111,W02121,W02201,W02211,W02221;
wire W02002,W02012,W02022,W02102,W02112,W02122,W02202,W02212,W02222;
wire signed [4:0] c00000,c01000,c02000;
wire signed [4:0] c00010,c01010,c02010;
wire signed [4:0] c00020,c01020,c02020;
wire signed [4:0] c00030,c01030,c02030;
wire signed [4:0] c00040,c01040,c02040;
wire signed [4:0] c00050,c01050,c02050;
wire signed [4:0] c00060,c01060,c02060;
wire signed [4:0] c00070,c01070,c02070;
wire signed [4:0] c00080,c01080,c02080;
wire signed [4:0] c00090,c01090,c02090;
wire signed [4:0] c000A0,c010A0,c020A0;
wire signed [4:0] c000B0,c010B0,c020B0;
wire signed [4:0] c000C0,c010C0,c020C0;
wire signed [4:0] c000D0,c010D0,c020D0;
wire signed [4:0] c00100,c01100,c02100;
wire signed [4:0] c00110,c01110,c02110;
wire signed [4:0] c00120,c01120,c02120;
wire signed [4:0] c00130,c01130,c02130;
wire signed [4:0] c00140,c01140,c02140;
wire signed [4:0] c00150,c01150,c02150;
wire signed [4:0] c00160,c01160,c02160;
wire signed [4:0] c00170,c01170,c02170;
wire signed [4:0] c00180,c01180,c02180;
wire signed [4:0] c00190,c01190,c02190;
wire signed [4:0] c001A0,c011A0,c021A0;
wire signed [4:0] c001B0,c011B0,c021B0;
wire signed [4:0] c001C0,c011C0,c021C0;
wire signed [4:0] c001D0,c011D0,c021D0;
wire signed [4:0] c00200,c01200,c02200;
wire signed [4:0] c00210,c01210,c02210;
wire signed [4:0] c00220,c01220,c02220;
wire signed [4:0] c00230,c01230,c02230;
wire signed [4:0] c00240,c01240,c02240;
wire signed [4:0] c00250,c01250,c02250;
wire signed [4:0] c00260,c01260,c02260;
wire signed [4:0] c00270,c01270,c02270;
wire signed [4:0] c00280,c01280,c02280;
wire signed [4:0] c00290,c01290,c02290;
wire signed [4:0] c002A0,c012A0,c022A0;
wire signed [4:0] c002B0,c012B0,c022B0;
wire signed [4:0] c002C0,c012C0,c022C0;
wire signed [4:0] c002D0,c012D0,c022D0;
wire signed [4:0] c00300,c01300,c02300;
wire signed [4:0] c00310,c01310,c02310;
wire signed [4:0] c00320,c01320,c02320;
wire signed [4:0] c00330,c01330,c02330;
wire signed [4:0] c00340,c01340,c02340;
wire signed [4:0] c00350,c01350,c02350;
wire signed [4:0] c00360,c01360,c02360;
wire signed [4:0] c00370,c01370,c02370;
wire signed [4:0] c00380,c01380,c02380;
wire signed [4:0] c00390,c01390,c02390;
wire signed [4:0] c003A0,c013A0,c023A0;
wire signed [4:0] c003B0,c013B0,c023B0;
wire signed [4:0] c003C0,c013C0,c023C0;
wire signed [4:0] c003D0,c013D0,c023D0;
wire signed [4:0] c00400,c01400,c02400;
wire signed [4:0] c00410,c01410,c02410;
wire signed [4:0] c00420,c01420,c02420;
wire signed [4:0] c00430,c01430,c02430;
wire signed [4:0] c00440,c01440,c02440;
wire signed [4:0] c00450,c01450,c02450;
wire signed [4:0] c00460,c01460,c02460;
wire signed [4:0] c00470,c01470,c02470;
wire signed [4:0] c00480,c01480,c02480;
wire signed [4:0] c00490,c01490,c02490;
wire signed [4:0] c004A0,c014A0,c024A0;
wire signed [4:0] c004B0,c014B0,c024B0;
wire signed [4:0] c004C0,c014C0,c024C0;
wire signed [4:0] c004D0,c014D0,c024D0;
wire signed [4:0] c00500,c01500,c02500;
wire signed [4:0] c00510,c01510,c02510;
wire signed [4:0] c00520,c01520,c02520;
wire signed [4:0] c00530,c01530,c02530;
wire signed [4:0] c00540,c01540,c02540;
wire signed [4:0] c00550,c01550,c02550;
wire signed [4:0] c00560,c01560,c02560;
wire signed [4:0] c00570,c01570,c02570;
wire signed [4:0] c00580,c01580,c02580;
wire signed [4:0] c00590,c01590,c02590;
wire signed [4:0] c005A0,c015A0,c025A0;
wire signed [4:0] c005B0,c015B0,c025B0;
wire signed [4:0] c005C0,c015C0,c025C0;
wire signed [4:0] c005D0,c015D0,c025D0;
wire signed [4:0] c00600,c01600,c02600;
wire signed [4:0] c00610,c01610,c02610;
wire signed [4:0] c00620,c01620,c02620;
wire signed [4:0] c00630,c01630,c02630;
wire signed [4:0] c00640,c01640,c02640;
wire signed [4:0] c00650,c01650,c02650;
wire signed [4:0] c00660,c01660,c02660;
wire signed [4:0] c00670,c01670,c02670;
wire signed [4:0] c00680,c01680,c02680;
wire signed [4:0] c00690,c01690,c02690;
wire signed [4:0] c006A0,c016A0,c026A0;
wire signed [4:0] c006B0,c016B0,c026B0;
wire signed [4:0] c006C0,c016C0,c026C0;
wire signed [4:0] c006D0,c016D0,c026D0;
wire signed [4:0] c00700,c01700,c02700;
wire signed [4:0] c00710,c01710,c02710;
wire signed [4:0] c00720,c01720,c02720;
wire signed [4:0] c00730,c01730,c02730;
wire signed [4:0] c00740,c01740,c02740;
wire signed [4:0] c00750,c01750,c02750;
wire signed [4:0] c00760,c01760,c02760;
wire signed [4:0] c00770,c01770,c02770;
wire signed [4:0] c00780,c01780,c02780;
wire signed [4:0] c00790,c01790,c02790;
wire signed [4:0] c007A0,c017A0,c027A0;
wire signed [4:0] c007B0,c017B0,c027B0;
wire signed [4:0] c007C0,c017C0,c027C0;
wire signed [4:0] c007D0,c017D0,c027D0;
wire signed [4:0] c00800,c01800,c02800;
wire signed [4:0] c00810,c01810,c02810;
wire signed [4:0] c00820,c01820,c02820;
wire signed [4:0] c00830,c01830,c02830;
wire signed [4:0] c00840,c01840,c02840;
wire signed [4:0] c00850,c01850,c02850;
wire signed [4:0] c00860,c01860,c02860;
wire signed [4:0] c00870,c01870,c02870;
wire signed [4:0] c00880,c01880,c02880;
wire signed [4:0] c00890,c01890,c02890;
wire signed [4:0] c008A0,c018A0,c028A0;
wire signed [4:0] c008B0,c018B0,c028B0;
wire signed [4:0] c008C0,c018C0,c028C0;
wire signed [4:0] c008D0,c018D0,c028D0;
wire signed [4:0] c00900,c01900,c02900;
wire signed [4:0] c00910,c01910,c02910;
wire signed [4:0] c00920,c01920,c02920;
wire signed [4:0] c00930,c01930,c02930;
wire signed [4:0] c00940,c01940,c02940;
wire signed [4:0] c00950,c01950,c02950;
wire signed [4:0] c00960,c01960,c02960;
wire signed [4:0] c00970,c01970,c02970;
wire signed [4:0] c00980,c01980,c02980;
wire signed [4:0] c00990,c01990,c02990;
wire signed [4:0] c009A0,c019A0,c029A0;
wire signed [4:0] c009B0,c019B0,c029B0;
wire signed [4:0] c009C0,c019C0,c029C0;
wire signed [4:0] c009D0,c019D0,c029D0;
wire signed [4:0] c00A00,c01A00,c02A00;
wire signed [4:0] c00A10,c01A10,c02A10;
wire signed [4:0] c00A20,c01A20,c02A20;
wire signed [4:0] c00A30,c01A30,c02A30;
wire signed [4:0] c00A40,c01A40,c02A40;
wire signed [4:0] c00A50,c01A50,c02A50;
wire signed [4:0] c00A60,c01A60,c02A60;
wire signed [4:0] c00A70,c01A70,c02A70;
wire signed [4:0] c00A80,c01A80,c02A80;
wire signed [4:0] c00A90,c01A90,c02A90;
wire signed [4:0] c00AA0,c01AA0,c02AA0;
wire signed [4:0] c00AB0,c01AB0,c02AB0;
wire signed [4:0] c00AC0,c01AC0,c02AC0;
wire signed [4:0] c00AD0,c01AD0,c02AD0;
wire signed [4:0] c00B00,c01B00,c02B00;
wire signed [4:0] c00B10,c01B10,c02B10;
wire signed [4:0] c00B20,c01B20,c02B20;
wire signed [4:0] c00B30,c01B30,c02B30;
wire signed [4:0] c00B40,c01B40,c02B40;
wire signed [4:0] c00B50,c01B50,c02B50;
wire signed [4:0] c00B60,c01B60,c02B60;
wire signed [4:0] c00B70,c01B70,c02B70;
wire signed [4:0] c00B80,c01B80,c02B80;
wire signed [4:0] c00B90,c01B90,c02B90;
wire signed [4:0] c00BA0,c01BA0,c02BA0;
wire signed [4:0] c00BB0,c01BB0,c02BB0;
wire signed [4:0] c00BC0,c01BC0,c02BC0;
wire signed [4:0] c00BD0,c01BD0,c02BD0;
wire signed [4:0] c00C00,c01C00,c02C00;
wire signed [4:0] c00C10,c01C10,c02C10;
wire signed [4:0] c00C20,c01C20,c02C20;
wire signed [4:0] c00C30,c01C30,c02C30;
wire signed [4:0] c00C40,c01C40,c02C40;
wire signed [4:0] c00C50,c01C50,c02C50;
wire signed [4:0] c00C60,c01C60,c02C60;
wire signed [4:0] c00C70,c01C70,c02C70;
wire signed [4:0] c00C80,c01C80,c02C80;
wire signed [4:0] c00C90,c01C90,c02C90;
wire signed [4:0] c00CA0,c01CA0,c02CA0;
wire signed [4:0] c00CB0,c01CB0,c02CB0;
wire signed [4:0] c00CC0,c01CC0,c02CC0;
wire signed [4:0] c00CD0,c01CD0,c02CD0;
wire signed [4:0] c00D00,c01D00,c02D00;
wire signed [4:0] c00D10,c01D10,c02D10;
wire signed [4:0] c00D20,c01D20,c02D20;
wire signed [4:0] c00D30,c01D30,c02D30;
wire signed [4:0] c00D40,c01D40,c02D40;
wire signed [4:0] c00D50,c01D50,c02D50;
wire signed [4:0] c00D60,c01D60,c02D60;
wire signed [4:0] c00D70,c01D70,c02D70;
wire signed [4:0] c00D80,c01D80,c02D80;
wire signed [4:0] c00D90,c01D90,c02D90;
wire signed [4:0] c00DA0,c01DA0,c02DA0;
wire signed [4:0] c00DB0,c01DB0,c02DB0;
wire signed [4:0] c00DC0,c01DC0,c02DC0;
wire signed [4:0] c00DD0,c01DD0,c02DD0;
wire signed [4:0] c00001,c01001,c02001;
wire signed [4:0] c00011,c01011,c02011;
wire signed [4:0] c00021,c01021,c02021;
wire signed [4:0] c00031,c01031,c02031;
wire signed [4:0] c00041,c01041,c02041;
wire signed [4:0] c00051,c01051,c02051;
wire signed [4:0] c00061,c01061,c02061;
wire signed [4:0] c00071,c01071,c02071;
wire signed [4:0] c00081,c01081,c02081;
wire signed [4:0] c00091,c01091,c02091;
wire signed [4:0] c000A1,c010A1,c020A1;
wire signed [4:0] c000B1,c010B1,c020B1;
wire signed [4:0] c000C1,c010C1,c020C1;
wire signed [4:0] c000D1,c010D1,c020D1;
wire signed [4:0] c00101,c01101,c02101;
wire signed [4:0] c00111,c01111,c02111;
wire signed [4:0] c00121,c01121,c02121;
wire signed [4:0] c00131,c01131,c02131;
wire signed [4:0] c00141,c01141,c02141;
wire signed [4:0] c00151,c01151,c02151;
wire signed [4:0] c00161,c01161,c02161;
wire signed [4:0] c00171,c01171,c02171;
wire signed [4:0] c00181,c01181,c02181;
wire signed [4:0] c00191,c01191,c02191;
wire signed [4:0] c001A1,c011A1,c021A1;
wire signed [4:0] c001B1,c011B1,c021B1;
wire signed [4:0] c001C1,c011C1,c021C1;
wire signed [4:0] c001D1,c011D1,c021D1;
wire signed [4:0] c00201,c01201,c02201;
wire signed [4:0] c00211,c01211,c02211;
wire signed [4:0] c00221,c01221,c02221;
wire signed [4:0] c00231,c01231,c02231;
wire signed [4:0] c00241,c01241,c02241;
wire signed [4:0] c00251,c01251,c02251;
wire signed [4:0] c00261,c01261,c02261;
wire signed [4:0] c00271,c01271,c02271;
wire signed [4:0] c00281,c01281,c02281;
wire signed [4:0] c00291,c01291,c02291;
wire signed [4:0] c002A1,c012A1,c022A1;
wire signed [4:0] c002B1,c012B1,c022B1;
wire signed [4:0] c002C1,c012C1,c022C1;
wire signed [4:0] c002D1,c012D1,c022D1;
wire signed [4:0] c00301,c01301,c02301;
wire signed [4:0] c00311,c01311,c02311;
wire signed [4:0] c00321,c01321,c02321;
wire signed [4:0] c00331,c01331,c02331;
wire signed [4:0] c00341,c01341,c02341;
wire signed [4:0] c00351,c01351,c02351;
wire signed [4:0] c00361,c01361,c02361;
wire signed [4:0] c00371,c01371,c02371;
wire signed [4:0] c00381,c01381,c02381;
wire signed [4:0] c00391,c01391,c02391;
wire signed [4:0] c003A1,c013A1,c023A1;
wire signed [4:0] c003B1,c013B1,c023B1;
wire signed [4:0] c003C1,c013C1,c023C1;
wire signed [4:0] c003D1,c013D1,c023D1;
wire signed [4:0] c00401,c01401,c02401;
wire signed [4:0] c00411,c01411,c02411;
wire signed [4:0] c00421,c01421,c02421;
wire signed [4:0] c00431,c01431,c02431;
wire signed [4:0] c00441,c01441,c02441;
wire signed [4:0] c00451,c01451,c02451;
wire signed [4:0] c00461,c01461,c02461;
wire signed [4:0] c00471,c01471,c02471;
wire signed [4:0] c00481,c01481,c02481;
wire signed [4:0] c00491,c01491,c02491;
wire signed [4:0] c004A1,c014A1,c024A1;
wire signed [4:0] c004B1,c014B1,c024B1;
wire signed [4:0] c004C1,c014C1,c024C1;
wire signed [4:0] c004D1,c014D1,c024D1;
wire signed [4:0] c00501,c01501,c02501;
wire signed [4:0] c00511,c01511,c02511;
wire signed [4:0] c00521,c01521,c02521;
wire signed [4:0] c00531,c01531,c02531;
wire signed [4:0] c00541,c01541,c02541;
wire signed [4:0] c00551,c01551,c02551;
wire signed [4:0] c00561,c01561,c02561;
wire signed [4:0] c00571,c01571,c02571;
wire signed [4:0] c00581,c01581,c02581;
wire signed [4:0] c00591,c01591,c02591;
wire signed [4:0] c005A1,c015A1,c025A1;
wire signed [4:0] c005B1,c015B1,c025B1;
wire signed [4:0] c005C1,c015C1,c025C1;
wire signed [4:0] c005D1,c015D1,c025D1;
wire signed [4:0] c00601,c01601,c02601;
wire signed [4:0] c00611,c01611,c02611;
wire signed [4:0] c00621,c01621,c02621;
wire signed [4:0] c00631,c01631,c02631;
wire signed [4:0] c00641,c01641,c02641;
wire signed [4:0] c00651,c01651,c02651;
wire signed [4:0] c00661,c01661,c02661;
wire signed [4:0] c00671,c01671,c02671;
wire signed [4:0] c00681,c01681,c02681;
wire signed [4:0] c00691,c01691,c02691;
wire signed [4:0] c006A1,c016A1,c026A1;
wire signed [4:0] c006B1,c016B1,c026B1;
wire signed [4:0] c006C1,c016C1,c026C1;
wire signed [4:0] c006D1,c016D1,c026D1;
wire signed [4:0] c00701,c01701,c02701;
wire signed [4:0] c00711,c01711,c02711;
wire signed [4:0] c00721,c01721,c02721;
wire signed [4:0] c00731,c01731,c02731;
wire signed [4:0] c00741,c01741,c02741;
wire signed [4:0] c00751,c01751,c02751;
wire signed [4:0] c00761,c01761,c02761;
wire signed [4:0] c00771,c01771,c02771;
wire signed [4:0] c00781,c01781,c02781;
wire signed [4:0] c00791,c01791,c02791;
wire signed [4:0] c007A1,c017A1,c027A1;
wire signed [4:0] c007B1,c017B1,c027B1;
wire signed [4:0] c007C1,c017C1,c027C1;
wire signed [4:0] c007D1,c017D1,c027D1;
wire signed [4:0] c00801,c01801,c02801;
wire signed [4:0] c00811,c01811,c02811;
wire signed [4:0] c00821,c01821,c02821;
wire signed [4:0] c00831,c01831,c02831;
wire signed [4:0] c00841,c01841,c02841;
wire signed [4:0] c00851,c01851,c02851;
wire signed [4:0] c00861,c01861,c02861;
wire signed [4:0] c00871,c01871,c02871;
wire signed [4:0] c00881,c01881,c02881;
wire signed [4:0] c00891,c01891,c02891;
wire signed [4:0] c008A1,c018A1,c028A1;
wire signed [4:0] c008B1,c018B1,c028B1;
wire signed [4:0] c008C1,c018C1,c028C1;
wire signed [4:0] c008D1,c018D1,c028D1;
wire signed [4:0] c00901,c01901,c02901;
wire signed [4:0] c00911,c01911,c02911;
wire signed [4:0] c00921,c01921,c02921;
wire signed [4:0] c00931,c01931,c02931;
wire signed [4:0] c00941,c01941,c02941;
wire signed [4:0] c00951,c01951,c02951;
wire signed [4:0] c00961,c01961,c02961;
wire signed [4:0] c00971,c01971,c02971;
wire signed [4:0] c00981,c01981,c02981;
wire signed [4:0] c00991,c01991,c02991;
wire signed [4:0] c009A1,c019A1,c029A1;
wire signed [4:0] c009B1,c019B1,c029B1;
wire signed [4:0] c009C1,c019C1,c029C1;
wire signed [4:0] c009D1,c019D1,c029D1;
wire signed [4:0] c00A01,c01A01,c02A01;
wire signed [4:0] c00A11,c01A11,c02A11;
wire signed [4:0] c00A21,c01A21,c02A21;
wire signed [4:0] c00A31,c01A31,c02A31;
wire signed [4:0] c00A41,c01A41,c02A41;
wire signed [4:0] c00A51,c01A51,c02A51;
wire signed [4:0] c00A61,c01A61,c02A61;
wire signed [4:0] c00A71,c01A71,c02A71;
wire signed [4:0] c00A81,c01A81,c02A81;
wire signed [4:0] c00A91,c01A91,c02A91;
wire signed [4:0] c00AA1,c01AA1,c02AA1;
wire signed [4:0] c00AB1,c01AB1,c02AB1;
wire signed [4:0] c00AC1,c01AC1,c02AC1;
wire signed [4:0] c00AD1,c01AD1,c02AD1;
wire signed [4:0] c00B01,c01B01,c02B01;
wire signed [4:0] c00B11,c01B11,c02B11;
wire signed [4:0] c00B21,c01B21,c02B21;
wire signed [4:0] c00B31,c01B31,c02B31;
wire signed [4:0] c00B41,c01B41,c02B41;
wire signed [4:0] c00B51,c01B51,c02B51;
wire signed [4:0] c00B61,c01B61,c02B61;
wire signed [4:0] c00B71,c01B71,c02B71;
wire signed [4:0] c00B81,c01B81,c02B81;
wire signed [4:0] c00B91,c01B91,c02B91;
wire signed [4:0] c00BA1,c01BA1,c02BA1;
wire signed [4:0] c00BB1,c01BB1,c02BB1;
wire signed [4:0] c00BC1,c01BC1,c02BC1;
wire signed [4:0] c00BD1,c01BD1,c02BD1;
wire signed [4:0] c00C01,c01C01,c02C01;
wire signed [4:0] c00C11,c01C11,c02C11;
wire signed [4:0] c00C21,c01C21,c02C21;
wire signed [4:0] c00C31,c01C31,c02C31;
wire signed [4:0] c00C41,c01C41,c02C41;
wire signed [4:0] c00C51,c01C51,c02C51;
wire signed [4:0] c00C61,c01C61,c02C61;
wire signed [4:0] c00C71,c01C71,c02C71;
wire signed [4:0] c00C81,c01C81,c02C81;
wire signed [4:0] c00C91,c01C91,c02C91;
wire signed [4:0] c00CA1,c01CA1,c02CA1;
wire signed [4:0] c00CB1,c01CB1,c02CB1;
wire signed [4:0] c00CC1,c01CC1,c02CC1;
wire signed [4:0] c00CD1,c01CD1,c02CD1;
wire signed [4:0] c00D01,c01D01,c02D01;
wire signed [4:0] c00D11,c01D11,c02D11;
wire signed [4:0] c00D21,c01D21,c02D21;
wire signed [4:0] c00D31,c01D31,c02D31;
wire signed [4:0] c00D41,c01D41,c02D41;
wire signed [4:0] c00D51,c01D51,c02D51;
wire signed [4:0] c00D61,c01D61,c02D61;
wire signed [4:0] c00D71,c01D71,c02D71;
wire signed [4:0] c00D81,c01D81,c02D81;
wire signed [4:0] c00D91,c01D91,c02D91;
wire signed [4:0] c00DA1,c01DA1,c02DA1;
wire signed [4:0] c00DB1,c01DB1,c02DB1;
wire signed [4:0] c00DC1,c01DC1,c02DC1;
wire signed [4:0] c00DD1,c01DD1,c02DD1;
wire signed [4:0] c00002,c01002,c02002;
wire signed [4:0] c00012,c01012,c02012;
wire signed [4:0] c00022,c01022,c02022;
wire signed [4:0] c00032,c01032,c02032;
wire signed [4:0] c00042,c01042,c02042;
wire signed [4:0] c00052,c01052,c02052;
wire signed [4:0] c00062,c01062,c02062;
wire signed [4:0] c00072,c01072,c02072;
wire signed [4:0] c00082,c01082,c02082;
wire signed [4:0] c00092,c01092,c02092;
wire signed [4:0] c000A2,c010A2,c020A2;
wire signed [4:0] c000B2,c010B2,c020B2;
wire signed [4:0] c000C2,c010C2,c020C2;
wire signed [4:0] c000D2,c010D2,c020D2;
wire signed [4:0] c00102,c01102,c02102;
wire signed [4:0] c00112,c01112,c02112;
wire signed [4:0] c00122,c01122,c02122;
wire signed [4:0] c00132,c01132,c02132;
wire signed [4:0] c00142,c01142,c02142;
wire signed [4:0] c00152,c01152,c02152;
wire signed [4:0] c00162,c01162,c02162;
wire signed [4:0] c00172,c01172,c02172;
wire signed [4:0] c00182,c01182,c02182;
wire signed [4:0] c00192,c01192,c02192;
wire signed [4:0] c001A2,c011A2,c021A2;
wire signed [4:0] c001B2,c011B2,c021B2;
wire signed [4:0] c001C2,c011C2,c021C2;
wire signed [4:0] c001D2,c011D2,c021D2;
wire signed [4:0] c00202,c01202,c02202;
wire signed [4:0] c00212,c01212,c02212;
wire signed [4:0] c00222,c01222,c02222;
wire signed [4:0] c00232,c01232,c02232;
wire signed [4:0] c00242,c01242,c02242;
wire signed [4:0] c00252,c01252,c02252;
wire signed [4:0] c00262,c01262,c02262;
wire signed [4:0] c00272,c01272,c02272;
wire signed [4:0] c00282,c01282,c02282;
wire signed [4:0] c00292,c01292,c02292;
wire signed [4:0] c002A2,c012A2,c022A2;
wire signed [4:0] c002B2,c012B2,c022B2;
wire signed [4:0] c002C2,c012C2,c022C2;
wire signed [4:0] c002D2,c012D2,c022D2;
wire signed [4:0] c00302,c01302,c02302;
wire signed [4:0] c00312,c01312,c02312;
wire signed [4:0] c00322,c01322,c02322;
wire signed [4:0] c00332,c01332,c02332;
wire signed [4:0] c00342,c01342,c02342;
wire signed [4:0] c00352,c01352,c02352;
wire signed [4:0] c00362,c01362,c02362;
wire signed [4:0] c00372,c01372,c02372;
wire signed [4:0] c00382,c01382,c02382;
wire signed [4:0] c00392,c01392,c02392;
wire signed [4:0] c003A2,c013A2,c023A2;
wire signed [4:0] c003B2,c013B2,c023B2;
wire signed [4:0] c003C2,c013C2,c023C2;
wire signed [4:0] c003D2,c013D2,c023D2;
wire signed [4:0] c00402,c01402,c02402;
wire signed [4:0] c00412,c01412,c02412;
wire signed [4:0] c00422,c01422,c02422;
wire signed [4:0] c00432,c01432,c02432;
wire signed [4:0] c00442,c01442,c02442;
wire signed [4:0] c00452,c01452,c02452;
wire signed [4:0] c00462,c01462,c02462;
wire signed [4:0] c00472,c01472,c02472;
wire signed [4:0] c00482,c01482,c02482;
wire signed [4:0] c00492,c01492,c02492;
wire signed [4:0] c004A2,c014A2,c024A2;
wire signed [4:0] c004B2,c014B2,c024B2;
wire signed [4:0] c004C2,c014C2,c024C2;
wire signed [4:0] c004D2,c014D2,c024D2;
wire signed [4:0] c00502,c01502,c02502;
wire signed [4:0] c00512,c01512,c02512;
wire signed [4:0] c00522,c01522,c02522;
wire signed [4:0] c00532,c01532,c02532;
wire signed [4:0] c00542,c01542,c02542;
wire signed [4:0] c00552,c01552,c02552;
wire signed [4:0] c00562,c01562,c02562;
wire signed [4:0] c00572,c01572,c02572;
wire signed [4:0] c00582,c01582,c02582;
wire signed [4:0] c00592,c01592,c02592;
wire signed [4:0] c005A2,c015A2,c025A2;
wire signed [4:0] c005B2,c015B2,c025B2;
wire signed [4:0] c005C2,c015C2,c025C2;
wire signed [4:0] c005D2,c015D2,c025D2;
wire signed [4:0] c00602,c01602,c02602;
wire signed [4:0] c00612,c01612,c02612;
wire signed [4:0] c00622,c01622,c02622;
wire signed [4:0] c00632,c01632,c02632;
wire signed [4:0] c00642,c01642,c02642;
wire signed [4:0] c00652,c01652,c02652;
wire signed [4:0] c00662,c01662,c02662;
wire signed [4:0] c00672,c01672,c02672;
wire signed [4:0] c00682,c01682,c02682;
wire signed [4:0] c00692,c01692,c02692;
wire signed [4:0] c006A2,c016A2,c026A2;
wire signed [4:0] c006B2,c016B2,c026B2;
wire signed [4:0] c006C2,c016C2,c026C2;
wire signed [4:0] c006D2,c016D2,c026D2;
wire signed [4:0] c00702,c01702,c02702;
wire signed [4:0] c00712,c01712,c02712;
wire signed [4:0] c00722,c01722,c02722;
wire signed [4:0] c00732,c01732,c02732;
wire signed [4:0] c00742,c01742,c02742;
wire signed [4:0] c00752,c01752,c02752;
wire signed [4:0] c00762,c01762,c02762;
wire signed [4:0] c00772,c01772,c02772;
wire signed [4:0] c00782,c01782,c02782;
wire signed [4:0] c00792,c01792,c02792;
wire signed [4:0] c007A2,c017A2,c027A2;
wire signed [4:0] c007B2,c017B2,c027B2;
wire signed [4:0] c007C2,c017C2,c027C2;
wire signed [4:0] c007D2,c017D2,c027D2;
wire signed [4:0] c00802,c01802,c02802;
wire signed [4:0] c00812,c01812,c02812;
wire signed [4:0] c00822,c01822,c02822;
wire signed [4:0] c00832,c01832,c02832;
wire signed [4:0] c00842,c01842,c02842;
wire signed [4:0] c00852,c01852,c02852;
wire signed [4:0] c00862,c01862,c02862;
wire signed [4:0] c00872,c01872,c02872;
wire signed [4:0] c00882,c01882,c02882;
wire signed [4:0] c00892,c01892,c02892;
wire signed [4:0] c008A2,c018A2,c028A2;
wire signed [4:0] c008B2,c018B2,c028B2;
wire signed [4:0] c008C2,c018C2,c028C2;
wire signed [4:0] c008D2,c018D2,c028D2;
wire signed [4:0] c00902,c01902,c02902;
wire signed [4:0] c00912,c01912,c02912;
wire signed [4:0] c00922,c01922,c02922;
wire signed [4:0] c00932,c01932,c02932;
wire signed [4:0] c00942,c01942,c02942;
wire signed [4:0] c00952,c01952,c02952;
wire signed [4:0] c00962,c01962,c02962;
wire signed [4:0] c00972,c01972,c02972;
wire signed [4:0] c00982,c01982,c02982;
wire signed [4:0] c00992,c01992,c02992;
wire signed [4:0] c009A2,c019A2,c029A2;
wire signed [4:0] c009B2,c019B2,c029B2;
wire signed [4:0] c009C2,c019C2,c029C2;
wire signed [4:0] c009D2,c019D2,c029D2;
wire signed [4:0] c00A02,c01A02,c02A02;
wire signed [4:0] c00A12,c01A12,c02A12;
wire signed [4:0] c00A22,c01A22,c02A22;
wire signed [4:0] c00A32,c01A32,c02A32;
wire signed [4:0] c00A42,c01A42,c02A42;
wire signed [4:0] c00A52,c01A52,c02A52;
wire signed [4:0] c00A62,c01A62,c02A62;
wire signed [4:0] c00A72,c01A72,c02A72;
wire signed [4:0] c00A82,c01A82,c02A82;
wire signed [4:0] c00A92,c01A92,c02A92;
wire signed [4:0] c00AA2,c01AA2,c02AA2;
wire signed [4:0] c00AB2,c01AB2,c02AB2;
wire signed [4:0] c00AC2,c01AC2,c02AC2;
wire signed [4:0] c00AD2,c01AD2,c02AD2;
wire signed [4:0] c00B02,c01B02,c02B02;
wire signed [4:0] c00B12,c01B12,c02B12;
wire signed [4:0] c00B22,c01B22,c02B22;
wire signed [4:0] c00B32,c01B32,c02B32;
wire signed [4:0] c00B42,c01B42,c02B42;
wire signed [4:0] c00B52,c01B52,c02B52;
wire signed [4:0] c00B62,c01B62,c02B62;
wire signed [4:0] c00B72,c01B72,c02B72;
wire signed [4:0] c00B82,c01B82,c02B82;
wire signed [4:0] c00B92,c01B92,c02B92;
wire signed [4:0] c00BA2,c01BA2,c02BA2;
wire signed [4:0] c00BB2,c01BB2,c02BB2;
wire signed [4:0] c00BC2,c01BC2,c02BC2;
wire signed [4:0] c00BD2,c01BD2,c02BD2;
wire signed [4:0] c00C02,c01C02,c02C02;
wire signed [4:0] c00C12,c01C12,c02C12;
wire signed [4:0] c00C22,c01C22,c02C22;
wire signed [4:0] c00C32,c01C32,c02C32;
wire signed [4:0] c00C42,c01C42,c02C42;
wire signed [4:0] c00C52,c01C52,c02C52;
wire signed [4:0] c00C62,c01C62,c02C62;
wire signed [4:0] c00C72,c01C72,c02C72;
wire signed [4:0] c00C82,c01C82,c02C82;
wire signed [4:0] c00C92,c01C92,c02C92;
wire signed [4:0] c00CA2,c01CA2,c02CA2;
wire signed [4:0] c00CB2,c01CB2,c02CB2;
wire signed [4:0] c00CC2,c01CC2,c02CC2;
wire signed [4:0] c00CD2,c01CD2,c02CD2;
wire signed [4:0] c00D02,c01D02,c02D02;
wire signed [4:0] c00D12,c01D12,c02D12;
wire signed [4:0] c00D22,c01D22,c02D22;
wire signed [4:0] c00D32,c01D32,c02D32;
wire signed [4:0] c00D42,c01D42,c02D42;
wire signed [4:0] c00D52,c01D52,c02D52;
wire signed [4:0] c00D62,c01D62,c02D62;
wire signed [4:0] c00D72,c01D72,c02D72;
wire signed [4:0] c00D82,c01D82,c02D82;
wire signed [4:0] c00D92,c01D92,c02D92;
wire signed [4:0] c00DA2,c01DA2,c02DA2;
wire signed [4:0] c00DB2,c01DB2,c02DB2;
wire signed [4:0] c00DC2,c01DC2,c02DC2;
wire signed [4:0] c00DD2,c01DD2,c02DD2;
wire signed [6:0] C0000;
wire A0000;
wire signed [6:0] C0010;
wire A0010;
wire signed [6:0] C0020;
wire A0020;
wire signed [6:0] C0030;
wire A0030;
wire signed [6:0] C0040;
wire A0040;
wire signed [6:0] C0050;
wire A0050;
wire signed [6:0] C0060;
wire A0060;
wire signed [6:0] C0070;
wire A0070;
wire signed [6:0] C0080;
wire A0080;
wire signed [6:0] C0090;
wire A0090;
wire signed [6:0] C00A0;
wire A00A0;
wire signed [6:0] C00B0;
wire A00B0;
wire signed [6:0] C00C0;
wire A00C0;
wire signed [6:0] C00D0;
wire A00D0;
wire signed [6:0] C0100;
wire A0100;
wire signed [6:0] C0110;
wire A0110;
wire signed [6:0] C0120;
wire A0120;
wire signed [6:0] C0130;
wire A0130;
wire signed [6:0] C0140;
wire A0140;
wire signed [6:0] C0150;
wire A0150;
wire signed [6:0] C0160;
wire A0160;
wire signed [6:0] C0170;
wire A0170;
wire signed [6:0] C0180;
wire A0180;
wire signed [6:0] C0190;
wire A0190;
wire signed [6:0] C01A0;
wire A01A0;
wire signed [6:0] C01B0;
wire A01B0;
wire signed [6:0] C01C0;
wire A01C0;
wire signed [6:0] C01D0;
wire A01D0;
wire signed [6:0] C0200;
wire A0200;
wire signed [6:0] C0210;
wire A0210;
wire signed [6:0] C0220;
wire A0220;
wire signed [6:0] C0230;
wire A0230;
wire signed [6:0] C0240;
wire A0240;
wire signed [6:0] C0250;
wire A0250;
wire signed [6:0] C0260;
wire A0260;
wire signed [6:0] C0270;
wire A0270;
wire signed [6:0] C0280;
wire A0280;
wire signed [6:0] C0290;
wire A0290;
wire signed [6:0] C02A0;
wire A02A0;
wire signed [6:0] C02B0;
wire A02B0;
wire signed [6:0] C02C0;
wire A02C0;
wire signed [6:0] C02D0;
wire A02D0;
wire signed [6:0] C0300;
wire A0300;
wire signed [6:0] C0310;
wire A0310;
wire signed [6:0] C0320;
wire A0320;
wire signed [6:0] C0330;
wire A0330;
wire signed [6:0] C0340;
wire A0340;
wire signed [6:0] C0350;
wire A0350;
wire signed [6:0] C0360;
wire A0360;
wire signed [6:0] C0370;
wire A0370;
wire signed [6:0] C0380;
wire A0380;
wire signed [6:0] C0390;
wire A0390;
wire signed [6:0] C03A0;
wire A03A0;
wire signed [6:0] C03B0;
wire A03B0;
wire signed [6:0] C03C0;
wire A03C0;
wire signed [6:0] C03D0;
wire A03D0;
wire signed [6:0] C0400;
wire A0400;
wire signed [6:0] C0410;
wire A0410;
wire signed [6:0] C0420;
wire A0420;
wire signed [6:0] C0430;
wire A0430;
wire signed [6:0] C0440;
wire A0440;
wire signed [6:0] C0450;
wire A0450;
wire signed [6:0] C0460;
wire A0460;
wire signed [6:0] C0470;
wire A0470;
wire signed [6:0] C0480;
wire A0480;
wire signed [6:0] C0490;
wire A0490;
wire signed [6:0] C04A0;
wire A04A0;
wire signed [6:0] C04B0;
wire A04B0;
wire signed [6:0] C04C0;
wire A04C0;
wire signed [6:0] C04D0;
wire A04D0;
wire signed [6:0] C0500;
wire A0500;
wire signed [6:0] C0510;
wire A0510;
wire signed [6:0] C0520;
wire A0520;
wire signed [6:0] C0530;
wire A0530;
wire signed [6:0] C0540;
wire A0540;
wire signed [6:0] C0550;
wire A0550;
wire signed [6:0] C0560;
wire A0560;
wire signed [6:0] C0570;
wire A0570;
wire signed [6:0] C0580;
wire A0580;
wire signed [6:0] C0590;
wire A0590;
wire signed [6:0] C05A0;
wire A05A0;
wire signed [6:0] C05B0;
wire A05B0;
wire signed [6:0] C05C0;
wire A05C0;
wire signed [6:0] C05D0;
wire A05D0;
wire signed [6:0] C0600;
wire A0600;
wire signed [6:0] C0610;
wire A0610;
wire signed [6:0] C0620;
wire A0620;
wire signed [6:0] C0630;
wire A0630;
wire signed [6:0] C0640;
wire A0640;
wire signed [6:0] C0650;
wire A0650;
wire signed [6:0] C0660;
wire A0660;
wire signed [6:0] C0670;
wire A0670;
wire signed [6:0] C0680;
wire A0680;
wire signed [6:0] C0690;
wire A0690;
wire signed [6:0] C06A0;
wire A06A0;
wire signed [6:0] C06B0;
wire A06B0;
wire signed [6:0] C06C0;
wire A06C0;
wire signed [6:0] C06D0;
wire A06D0;
wire signed [6:0] C0700;
wire A0700;
wire signed [6:0] C0710;
wire A0710;
wire signed [6:0] C0720;
wire A0720;
wire signed [6:0] C0730;
wire A0730;
wire signed [6:0] C0740;
wire A0740;
wire signed [6:0] C0750;
wire A0750;
wire signed [6:0] C0760;
wire A0760;
wire signed [6:0] C0770;
wire A0770;
wire signed [6:0] C0780;
wire A0780;
wire signed [6:0] C0790;
wire A0790;
wire signed [6:0] C07A0;
wire A07A0;
wire signed [6:0] C07B0;
wire A07B0;
wire signed [6:0] C07C0;
wire A07C0;
wire signed [6:0] C07D0;
wire A07D0;
wire signed [6:0] C0800;
wire A0800;
wire signed [6:0] C0810;
wire A0810;
wire signed [6:0] C0820;
wire A0820;
wire signed [6:0] C0830;
wire A0830;
wire signed [6:0] C0840;
wire A0840;
wire signed [6:0] C0850;
wire A0850;
wire signed [6:0] C0860;
wire A0860;
wire signed [6:0] C0870;
wire A0870;
wire signed [6:0] C0880;
wire A0880;
wire signed [6:0] C0890;
wire A0890;
wire signed [6:0] C08A0;
wire A08A0;
wire signed [6:0] C08B0;
wire A08B0;
wire signed [6:0] C08C0;
wire A08C0;
wire signed [6:0] C08D0;
wire A08D0;
wire signed [6:0] C0900;
wire A0900;
wire signed [6:0] C0910;
wire A0910;
wire signed [6:0] C0920;
wire A0920;
wire signed [6:0] C0930;
wire A0930;
wire signed [6:0] C0940;
wire A0940;
wire signed [6:0] C0950;
wire A0950;
wire signed [6:0] C0960;
wire A0960;
wire signed [6:0] C0970;
wire A0970;
wire signed [6:0] C0980;
wire A0980;
wire signed [6:0] C0990;
wire A0990;
wire signed [6:0] C09A0;
wire A09A0;
wire signed [6:0] C09B0;
wire A09B0;
wire signed [6:0] C09C0;
wire A09C0;
wire signed [6:0] C09D0;
wire A09D0;
wire signed [6:0] C0A00;
wire A0A00;
wire signed [6:0] C0A10;
wire A0A10;
wire signed [6:0] C0A20;
wire A0A20;
wire signed [6:0] C0A30;
wire A0A30;
wire signed [6:0] C0A40;
wire A0A40;
wire signed [6:0] C0A50;
wire A0A50;
wire signed [6:0] C0A60;
wire A0A60;
wire signed [6:0] C0A70;
wire A0A70;
wire signed [6:0] C0A80;
wire A0A80;
wire signed [6:0] C0A90;
wire A0A90;
wire signed [6:0] C0AA0;
wire A0AA0;
wire signed [6:0] C0AB0;
wire A0AB0;
wire signed [6:0] C0AC0;
wire A0AC0;
wire signed [6:0] C0AD0;
wire A0AD0;
wire signed [6:0] C0B00;
wire A0B00;
wire signed [6:0] C0B10;
wire A0B10;
wire signed [6:0] C0B20;
wire A0B20;
wire signed [6:0] C0B30;
wire A0B30;
wire signed [6:0] C0B40;
wire A0B40;
wire signed [6:0] C0B50;
wire A0B50;
wire signed [6:0] C0B60;
wire A0B60;
wire signed [6:0] C0B70;
wire A0B70;
wire signed [6:0] C0B80;
wire A0B80;
wire signed [6:0] C0B90;
wire A0B90;
wire signed [6:0] C0BA0;
wire A0BA0;
wire signed [6:0] C0BB0;
wire A0BB0;
wire signed [6:0] C0BC0;
wire A0BC0;
wire signed [6:0] C0BD0;
wire A0BD0;
wire signed [6:0] C0C00;
wire A0C00;
wire signed [6:0] C0C10;
wire A0C10;
wire signed [6:0] C0C20;
wire A0C20;
wire signed [6:0] C0C30;
wire A0C30;
wire signed [6:0] C0C40;
wire A0C40;
wire signed [6:0] C0C50;
wire A0C50;
wire signed [6:0] C0C60;
wire A0C60;
wire signed [6:0] C0C70;
wire A0C70;
wire signed [6:0] C0C80;
wire A0C80;
wire signed [6:0] C0C90;
wire A0C90;
wire signed [6:0] C0CA0;
wire A0CA0;
wire signed [6:0] C0CB0;
wire A0CB0;
wire signed [6:0] C0CC0;
wire A0CC0;
wire signed [6:0] C0CD0;
wire A0CD0;
wire signed [6:0] C0D00;
wire A0D00;
wire signed [6:0] C0D10;
wire A0D10;
wire signed [6:0] C0D20;
wire A0D20;
wire signed [6:0] C0D30;
wire A0D30;
wire signed [6:0] C0D40;
wire A0D40;
wire signed [6:0] C0D50;
wire A0D50;
wire signed [6:0] C0D60;
wire A0D60;
wire signed [6:0] C0D70;
wire A0D70;
wire signed [6:0] C0D80;
wire A0D80;
wire signed [6:0] C0D90;
wire A0D90;
wire signed [6:0] C0DA0;
wire A0DA0;
wire signed [6:0] C0DB0;
wire A0DB0;
wire signed [6:0] C0DC0;
wire A0DC0;
wire signed [6:0] C0DD0;
wire A0DD0;
wire signed [6:0] C0001;
wire A0001;
wire signed [6:0] C0011;
wire A0011;
wire signed [6:0] C0021;
wire A0021;
wire signed [6:0] C0031;
wire A0031;
wire signed [6:0] C0041;
wire A0041;
wire signed [6:0] C0051;
wire A0051;
wire signed [6:0] C0061;
wire A0061;
wire signed [6:0] C0071;
wire A0071;
wire signed [6:0] C0081;
wire A0081;
wire signed [6:0] C0091;
wire A0091;
wire signed [6:0] C00A1;
wire A00A1;
wire signed [6:0] C00B1;
wire A00B1;
wire signed [6:0] C00C1;
wire A00C1;
wire signed [6:0] C00D1;
wire A00D1;
wire signed [6:0] C0101;
wire A0101;
wire signed [6:0] C0111;
wire A0111;
wire signed [6:0] C0121;
wire A0121;
wire signed [6:0] C0131;
wire A0131;
wire signed [6:0] C0141;
wire A0141;
wire signed [6:0] C0151;
wire A0151;
wire signed [6:0] C0161;
wire A0161;
wire signed [6:0] C0171;
wire A0171;
wire signed [6:0] C0181;
wire A0181;
wire signed [6:0] C0191;
wire A0191;
wire signed [6:0] C01A1;
wire A01A1;
wire signed [6:0] C01B1;
wire A01B1;
wire signed [6:0] C01C1;
wire A01C1;
wire signed [6:0] C01D1;
wire A01D1;
wire signed [6:0] C0201;
wire A0201;
wire signed [6:0] C0211;
wire A0211;
wire signed [6:0] C0221;
wire A0221;
wire signed [6:0] C0231;
wire A0231;
wire signed [6:0] C0241;
wire A0241;
wire signed [6:0] C0251;
wire A0251;
wire signed [6:0] C0261;
wire A0261;
wire signed [6:0] C0271;
wire A0271;
wire signed [6:0] C0281;
wire A0281;
wire signed [6:0] C0291;
wire A0291;
wire signed [6:0] C02A1;
wire A02A1;
wire signed [6:0] C02B1;
wire A02B1;
wire signed [6:0] C02C1;
wire A02C1;
wire signed [6:0] C02D1;
wire A02D1;
wire signed [6:0] C0301;
wire A0301;
wire signed [6:0] C0311;
wire A0311;
wire signed [6:0] C0321;
wire A0321;
wire signed [6:0] C0331;
wire A0331;
wire signed [6:0] C0341;
wire A0341;
wire signed [6:0] C0351;
wire A0351;
wire signed [6:0] C0361;
wire A0361;
wire signed [6:0] C0371;
wire A0371;
wire signed [6:0] C0381;
wire A0381;
wire signed [6:0] C0391;
wire A0391;
wire signed [6:0] C03A1;
wire A03A1;
wire signed [6:0] C03B1;
wire A03B1;
wire signed [6:0] C03C1;
wire A03C1;
wire signed [6:0] C03D1;
wire A03D1;
wire signed [6:0] C0401;
wire A0401;
wire signed [6:0] C0411;
wire A0411;
wire signed [6:0] C0421;
wire A0421;
wire signed [6:0] C0431;
wire A0431;
wire signed [6:0] C0441;
wire A0441;
wire signed [6:0] C0451;
wire A0451;
wire signed [6:0] C0461;
wire A0461;
wire signed [6:0] C0471;
wire A0471;
wire signed [6:0] C0481;
wire A0481;
wire signed [6:0] C0491;
wire A0491;
wire signed [6:0] C04A1;
wire A04A1;
wire signed [6:0] C04B1;
wire A04B1;
wire signed [6:0] C04C1;
wire A04C1;
wire signed [6:0] C04D1;
wire A04D1;
wire signed [6:0] C0501;
wire A0501;
wire signed [6:0] C0511;
wire A0511;
wire signed [6:0] C0521;
wire A0521;
wire signed [6:0] C0531;
wire A0531;
wire signed [6:0] C0541;
wire A0541;
wire signed [6:0] C0551;
wire A0551;
wire signed [6:0] C0561;
wire A0561;
wire signed [6:0] C0571;
wire A0571;
wire signed [6:0] C0581;
wire A0581;
wire signed [6:0] C0591;
wire A0591;
wire signed [6:0] C05A1;
wire A05A1;
wire signed [6:0] C05B1;
wire A05B1;
wire signed [6:0] C05C1;
wire A05C1;
wire signed [6:0] C05D1;
wire A05D1;
wire signed [6:0] C0601;
wire A0601;
wire signed [6:0] C0611;
wire A0611;
wire signed [6:0] C0621;
wire A0621;
wire signed [6:0] C0631;
wire A0631;
wire signed [6:0] C0641;
wire A0641;
wire signed [6:0] C0651;
wire A0651;
wire signed [6:0] C0661;
wire A0661;
wire signed [6:0] C0671;
wire A0671;
wire signed [6:0] C0681;
wire A0681;
wire signed [6:0] C0691;
wire A0691;
wire signed [6:0] C06A1;
wire A06A1;
wire signed [6:0] C06B1;
wire A06B1;
wire signed [6:0] C06C1;
wire A06C1;
wire signed [6:0] C06D1;
wire A06D1;
wire signed [6:0] C0701;
wire A0701;
wire signed [6:0] C0711;
wire A0711;
wire signed [6:0] C0721;
wire A0721;
wire signed [6:0] C0731;
wire A0731;
wire signed [6:0] C0741;
wire A0741;
wire signed [6:0] C0751;
wire A0751;
wire signed [6:0] C0761;
wire A0761;
wire signed [6:0] C0771;
wire A0771;
wire signed [6:0] C0781;
wire A0781;
wire signed [6:0] C0791;
wire A0791;
wire signed [6:0] C07A1;
wire A07A1;
wire signed [6:0] C07B1;
wire A07B1;
wire signed [6:0] C07C1;
wire A07C1;
wire signed [6:0] C07D1;
wire A07D1;
wire signed [6:0] C0801;
wire A0801;
wire signed [6:0] C0811;
wire A0811;
wire signed [6:0] C0821;
wire A0821;
wire signed [6:0] C0831;
wire A0831;
wire signed [6:0] C0841;
wire A0841;
wire signed [6:0] C0851;
wire A0851;
wire signed [6:0] C0861;
wire A0861;
wire signed [6:0] C0871;
wire A0871;
wire signed [6:0] C0881;
wire A0881;
wire signed [6:0] C0891;
wire A0891;
wire signed [6:0] C08A1;
wire A08A1;
wire signed [6:0] C08B1;
wire A08B1;
wire signed [6:0] C08C1;
wire A08C1;
wire signed [6:0] C08D1;
wire A08D1;
wire signed [6:0] C0901;
wire A0901;
wire signed [6:0] C0911;
wire A0911;
wire signed [6:0] C0921;
wire A0921;
wire signed [6:0] C0931;
wire A0931;
wire signed [6:0] C0941;
wire A0941;
wire signed [6:0] C0951;
wire A0951;
wire signed [6:0] C0961;
wire A0961;
wire signed [6:0] C0971;
wire A0971;
wire signed [6:0] C0981;
wire A0981;
wire signed [6:0] C0991;
wire A0991;
wire signed [6:0] C09A1;
wire A09A1;
wire signed [6:0] C09B1;
wire A09B1;
wire signed [6:0] C09C1;
wire A09C1;
wire signed [6:0] C09D1;
wire A09D1;
wire signed [6:0] C0A01;
wire A0A01;
wire signed [6:0] C0A11;
wire A0A11;
wire signed [6:0] C0A21;
wire A0A21;
wire signed [6:0] C0A31;
wire A0A31;
wire signed [6:0] C0A41;
wire A0A41;
wire signed [6:0] C0A51;
wire A0A51;
wire signed [6:0] C0A61;
wire A0A61;
wire signed [6:0] C0A71;
wire A0A71;
wire signed [6:0] C0A81;
wire A0A81;
wire signed [6:0] C0A91;
wire A0A91;
wire signed [6:0] C0AA1;
wire A0AA1;
wire signed [6:0] C0AB1;
wire A0AB1;
wire signed [6:0] C0AC1;
wire A0AC1;
wire signed [6:0] C0AD1;
wire A0AD1;
wire signed [6:0] C0B01;
wire A0B01;
wire signed [6:0] C0B11;
wire A0B11;
wire signed [6:0] C0B21;
wire A0B21;
wire signed [6:0] C0B31;
wire A0B31;
wire signed [6:0] C0B41;
wire A0B41;
wire signed [6:0] C0B51;
wire A0B51;
wire signed [6:0] C0B61;
wire A0B61;
wire signed [6:0] C0B71;
wire A0B71;
wire signed [6:0] C0B81;
wire A0B81;
wire signed [6:0] C0B91;
wire A0B91;
wire signed [6:0] C0BA1;
wire A0BA1;
wire signed [6:0] C0BB1;
wire A0BB1;
wire signed [6:0] C0BC1;
wire A0BC1;
wire signed [6:0] C0BD1;
wire A0BD1;
wire signed [6:0] C0C01;
wire A0C01;
wire signed [6:0] C0C11;
wire A0C11;
wire signed [6:0] C0C21;
wire A0C21;
wire signed [6:0] C0C31;
wire A0C31;
wire signed [6:0] C0C41;
wire A0C41;
wire signed [6:0] C0C51;
wire A0C51;
wire signed [6:0] C0C61;
wire A0C61;
wire signed [6:0] C0C71;
wire A0C71;
wire signed [6:0] C0C81;
wire A0C81;
wire signed [6:0] C0C91;
wire A0C91;
wire signed [6:0] C0CA1;
wire A0CA1;
wire signed [6:0] C0CB1;
wire A0CB1;
wire signed [6:0] C0CC1;
wire A0CC1;
wire signed [6:0] C0CD1;
wire A0CD1;
wire signed [6:0] C0D01;
wire A0D01;
wire signed [6:0] C0D11;
wire A0D11;
wire signed [6:0] C0D21;
wire A0D21;
wire signed [6:0] C0D31;
wire A0D31;
wire signed [6:0] C0D41;
wire A0D41;
wire signed [6:0] C0D51;
wire A0D51;
wire signed [6:0] C0D61;
wire A0D61;
wire signed [6:0] C0D71;
wire A0D71;
wire signed [6:0] C0D81;
wire A0D81;
wire signed [6:0] C0D91;
wire A0D91;
wire signed [6:0] C0DA1;
wire A0DA1;
wire signed [6:0] C0DB1;
wire A0DB1;
wire signed [6:0] C0DC1;
wire A0DC1;
wire signed [6:0] C0DD1;
wire A0DD1;
wire signed [6:0] C0002;
wire A0002;
wire signed [6:0] C0012;
wire A0012;
wire signed [6:0] C0022;
wire A0022;
wire signed [6:0] C0032;
wire A0032;
wire signed [6:0] C0042;
wire A0042;
wire signed [6:0] C0052;
wire A0052;
wire signed [6:0] C0062;
wire A0062;
wire signed [6:0] C0072;
wire A0072;
wire signed [6:0] C0082;
wire A0082;
wire signed [6:0] C0092;
wire A0092;
wire signed [6:0] C00A2;
wire A00A2;
wire signed [6:0] C00B2;
wire A00B2;
wire signed [6:0] C00C2;
wire A00C2;
wire signed [6:0] C00D2;
wire A00D2;
wire signed [6:0] C0102;
wire A0102;
wire signed [6:0] C0112;
wire A0112;
wire signed [6:0] C0122;
wire A0122;
wire signed [6:0] C0132;
wire A0132;
wire signed [6:0] C0142;
wire A0142;
wire signed [6:0] C0152;
wire A0152;
wire signed [6:0] C0162;
wire A0162;
wire signed [6:0] C0172;
wire A0172;
wire signed [6:0] C0182;
wire A0182;
wire signed [6:0] C0192;
wire A0192;
wire signed [6:0] C01A2;
wire A01A2;
wire signed [6:0] C01B2;
wire A01B2;
wire signed [6:0] C01C2;
wire A01C2;
wire signed [6:0] C01D2;
wire A01D2;
wire signed [6:0] C0202;
wire A0202;
wire signed [6:0] C0212;
wire A0212;
wire signed [6:0] C0222;
wire A0222;
wire signed [6:0] C0232;
wire A0232;
wire signed [6:0] C0242;
wire A0242;
wire signed [6:0] C0252;
wire A0252;
wire signed [6:0] C0262;
wire A0262;
wire signed [6:0] C0272;
wire A0272;
wire signed [6:0] C0282;
wire A0282;
wire signed [6:0] C0292;
wire A0292;
wire signed [6:0] C02A2;
wire A02A2;
wire signed [6:0] C02B2;
wire A02B2;
wire signed [6:0] C02C2;
wire A02C2;
wire signed [6:0] C02D2;
wire A02D2;
wire signed [6:0] C0302;
wire A0302;
wire signed [6:0] C0312;
wire A0312;
wire signed [6:0] C0322;
wire A0322;
wire signed [6:0] C0332;
wire A0332;
wire signed [6:0] C0342;
wire A0342;
wire signed [6:0] C0352;
wire A0352;
wire signed [6:0] C0362;
wire A0362;
wire signed [6:0] C0372;
wire A0372;
wire signed [6:0] C0382;
wire A0382;
wire signed [6:0] C0392;
wire A0392;
wire signed [6:0] C03A2;
wire A03A2;
wire signed [6:0] C03B2;
wire A03B2;
wire signed [6:0] C03C2;
wire A03C2;
wire signed [6:0] C03D2;
wire A03D2;
wire signed [6:0] C0402;
wire A0402;
wire signed [6:0] C0412;
wire A0412;
wire signed [6:0] C0422;
wire A0422;
wire signed [6:0] C0432;
wire A0432;
wire signed [6:0] C0442;
wire A0442;
wire signed [6:0] C0452;
wire A0452;
wire signed [6:0] C0462;
wire A0462;
wire signed [6:0] C0472;
wire A0472;
wire signed [6:0] C0482;
wire A0482;
wire signed [6:0] C0492;
wire A0492;
wire signed [6:0] C04A2;
wire A04A2;
wire signed [6:0] C04B2;
wire A04B2;
wire signed [6:0] C04C2;
wire A04C2;
wire signed [6:0] C04D2;
wire A04D2;
wire signed [6:0] C0502;
wire A0502;
wire signed [6:0] C0512;
wire A0512;
wire signed [6:0] C0522;
wire A0522;
wire signed [6:0] C0532;
wire A0532;
wire signed [6:0] C0542;
wire A0542;
wire signed [6:0] C0552;
wire A0552;
wire signed [6:0] C0562;
wire A0562;
wire signed [6:0] C0572;
wire A0572;
wire signed [6:0] C0582;
wire A0582;
wire signed [6:0] C0592;
wire A0592;
wire signed [6:0] C05A2;
wire A05A2;
wire signed [6:0] C05B2;
wire A05B2;
wire signed [6:0] C05C2;
wire A05C2;
wire signed [6:0] C05D2;
wire A05D2;
wire signed [6:0] C0602;
wire A0602;
wire signed [6:0] C0612;
wire A0612;
wire signed [6:0] C0622;
wire A0622;
wire signed [6:0] C0632;
wire A0632;
wire signed [6:0] C0642;
wire A0642;
wire signed [6:0] C0652;
wire A0652;
wire signed [6:0] C0662;
wire A0662;
wire signed [6:0] C0672;
wire A0672;
wire signed [6:0] C0682;
wire A0682;
wire signed [6:0] C0692;
wire A0692;
wire signed [6:0] C06A2;
wire A06A2;
wire signed [6:0] C06B2;
wire A06B2;
wire signed [6:0] C06C2;
wire A06C2;
wire signed [6:0] C06D2;
wire A06D2;
wire signed [6:0] C0702;
wire A0702;
wire signed [6:0] C0712;
wire A0712;
wire signed [6:0] C0722;
wire A0722;
wire signed [6:0] C0732;
wire A0732;
wire signed [6:0] C0742;
wire A0742;
wire signed [6:0] C0752;
wire A0752;
wire signed [6:0] C0762;
wire A0762;
wire signed [6:0] C0772;
wire A0772;
wire signed [6:0] C0782;
wire A0782;
wire signed [6:0] C0792;
wire A0792;
wire signed [6:0] C07A2;
wire A07A2;
wire signed [6:0] C07B2;
wire A07B2;
wire signed [6:0] C07C2;
wire A07C2;
wire signed [6:0] C07D2;
wire A07D2;
wire signed [6:0] C0802;
wire A0802;
wire signed [6:0] C0812;
wire A0812;
wire signed [6:0] C0822;
wire A0822;
wire signed [6:0] C0832;
wire A0832;
wire signed [6:0] C0842;
wire A0842;
wire signed [6:0] C0852;
wire A0852;
wire signed [6:0] C0862;
wire A0862;
wire signed [6:0] C0872;
wire A0872;
wire signed [6:0] C0882;
wire A0882;
wire signed [6:0] C0892;
wire A0892;
wire signed [6:0] C08A2;
wire A08A2;
wire signed [6:0] C08B2;
wire A08B2;
wire signed [6:0] C08C2;
wire A08C2;
wire signed [6:0] C08D2;
wire A08D2;
wire signed [6:0] C0902;
wire A0902;
wire signed [6:0] C0912;
wire A0912;
wire signed [6:0] C0922;
wire A0922;
wire signed [6:0] C0932;
wire A0932;
wire signed [6:0] C0942;
wire A0942;
wire signed [6:0] C0952;
wire A0952;
wire signed [6:0] C0962;
wire A0962;
wire signed [6:0] C0972;
wire A0972;
wire signed [6:0] C0982;
wire A0982;
wire signed [6:0] C0992;
wire A0992;
wire signed [6:0] C09A2;
wire A09A2;
wire signed [6:0] C09B2;
wire A09B2;
wire signed [6:0] C09C2;
wire A09C2;
wire signed [6:0] C09D2;
wire A09D2;
wire signed [6:0] C0A02;
wire A0A02;
wire signed [6:0] C0A12;
wire A0A12;
wire signed [6:0] C0A22;
wire A0A22;
wire signed [6:0] C0A32;
wire A0A32;
wire signed [6:0] C0A42;
wire A0A42;
wire signed [6:0] C0A52;
wire A0A52;
wire signed [6:0] C0A62;
wire A0A62;
wire signed [6:0] C0A72;
wire A0A72;
wire signed [6:0] C0A82;
wire A0A82;
wire signed [6:0] C0A92;
wire A0A92;
wire signed [6:0] C0AA2;
wire A0AA2;
wire signed [6:0] C0AB2;
wire A0AB2;
wire signed [6:0] C0AC2;
wire A0AC2;
wire signed [6:0] C0AD2;
wire A0AD2;
wire signed [6:0] C0B02;
wire A0B02;
wire signed [6:0] C0B12;
wire A0B12;
wire signed [6:0] C0B22;
wire A0B22;
wire signed [6:0] C0B32;
wire A0B32;
wire signed [6:0] C0B42;
wire A0B42;
wire signed [6:0] C0B52;
wire A0B52;
wire signed [6:0] C0B62;
wire A0B62;
wire signed [6:0] C0B72;
wire A0B72;
wire signed [6:0] C0B82;
wire A0B82;
wire signed [6:0] C0B92;
wire A0B92;
wire signed [6:0] C0BA2;
wire A0BA2;
wire signed [6:0] C0BB2;
wire A0BB2;
wire signed [6:0] C0BC2;
wire A0BC2;
wire signed [6:0] C0BD2;
wire A0BD2;
wire signed [6:0] C0C02;
wire A0C02;
wire signed [6:0] C0C12;
wire A0C12;
wire signed [6:0] C0C22;
wire A0C22;
wire signed [6:0] C0C32;
wire A0C32;
wire signed [6:0] C0C42;
wire A0C42;
wire signed [6:0] C0C52;
wire A0C52;
wire signed [6:0] C0C62;
wire A0C62;
wire signed [6:0] C0C72;
wire A0C72;
wire signed [6:0] C0C82;
wire A0C82;
wire signed [6:0] C0C92;
wire A0C92;
wire signed [6:0] C0CA2;
wire A0CA2;
wire signed [6:0] C0CB2;
wire A0CB2;
wire signed [6:0] C0CC2;
wire A0CC2;
wire signed [6:0] C0CD2;
wire A0CD2;
wire signed [6:0] C0D02;
wire A0D02;
wire signed [6:0] C0D12;
wire A0D12;
wire signed [6:0] C0D22;
wire A0D22;
wire signed [6:0] C0D32;
wire A0D32;
wire signed [6:0] C0D42;
wire A0D42;
wire signed [6:0] C0D52;
wire A0D52;
wire signed [6:0] C0D62;
wire A0D62;
wire signed [6:0] C0D72;
wire A0D72;
wire signed [6:0] C0D82;
wire A0D82;
wire signed [6:0] C0D92;
wire A0D92;
wire signed [6:0] C0DA2;
wire A0DA2;
wire signed [6:0] C0DB2;
wire A0DB2;
wire signed [6:0] C0DC2;
wire A0DC2;
wire signed [6:0] C0DD2;
wire A0DD2;
DFF_save_fm DFF_P0(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0000));
DFF_save_fm DFF_P1(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0010));
DFF_save_fm DFF_P2(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0020));
DFF_save_fm DFF_P3(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0030));
DFF_save_fm DFF_P4(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0040));
DFF_save_fm DFF_P5(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0050));
DFF_save_fm DFF_P6(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0060));
DFF_save_fm DFF_P7(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0070));
DFF_save_fm DFF_P8(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0080));
DFF_save_fm DFF_P9(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0090));
DFF_save_fm DFF_P10(.clk(clk),.rstn(rstn),.reset_value(1),.q(P00A0));
DFF_save_fm DFF_P11(.clk(clk),.rstn(rstn),.reset_value(1),.q(P00B0));
DFF_save_fm DFF_P12(.clk(clk),.rstn(rstn),.reset_value(1),.q(P00C0));
DFF_save_fm DFF_P13(.clk(clk),.rstn(rstn),.reset_value(1),.q(P00D0));
DFF_save_fm DFF_P14(.clk(clk),.rstn(rstn),.reset_value(1),.q(P00E0));
DFF_save_fm DFF_P15(.clk(clk),.rstn(rstn),.reset_value(1),.q(P00F0));
DFF_save_fm DFF_P16(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0100));
DFF_save_fm DFF_P17(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0110));
DFF_save_fm DFF_P18(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0120));
DFF_save_fm DFF_P19(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0130));
DFF_save_fm DFF_P20(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0140));
DFF_save_fm DFF_P21(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0150));
DFF_save_fm DFF_P22(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0160));
DFF_save_fm DFF_P23(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0170));
DFF_save_fm DFF_P24(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0180));
DFF_save_fm DFF_P25(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0190));
DFF_save_fm DFF_P26(.clk(clk),.rstn(rstn),.reset_value(1),.q(P01A0));
DFF_save_fm DFF_P27(.clk(clk),.rstn(rstn),.reset_value(0),.q(P01B0));
DFF_save_fm DFF_P28(.clk(clk),.rstn(rstn),.reset_value(0),.q(P01C0));
DFF_save_fm DFF_P29(.clk(clk),.rstn(rstn),.reset_value(1),.q(P01D0));
DFF_save_fm DFF_P30(.clk(clk),.rstn(rstn),.reset_value(1),.q(P01E0));
DFF_save_fm DFF_P31(.clk(clk),.rstn(rstn),.reset_value(1),.q(P01F0));
DFF_save_fm DFF_P32(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0200));
DFF_save_fm DFF_P33(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0210));
DFF_save_fm DFF_P34(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0220));
DFF_save_fm DFF_P35(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0230));
DFF_save_fm DFF_P36(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0240));
DFF_save_fm DFF_P37(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0250));
DFF_save_fm DFF_P38(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0260));
DFF_save_fm DFF_P39(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0270));
DFF_save_fm DFF_P40(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0280));
DFF_save_fm DFF_P41(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0290));
DFF_save_fm DFF_P42(.clk(clk),.rstn(rstn),.reset_value(1),.q(P02A0));
DFF_save_fm DFF_P43(.clk(clk),.rstn(rstn),.reset_value(0),.q(P02B0));
DFF_save_fm DFF_P44(.clk(clk),.rstn(rstn),.reset_value(0),.q(P02C0));
DFF_save_fm DFF_P45(.clk(clk),.rstn(rstn),.reset_value(1),.q(P02D0));
DFF_save_fm DFF_P46(.clk(clk),.rstn(rstn),.reset_value(1),.q(P02E0));
DFF_save_fm DFF_P47(.clk(clk),.rstn(rstn),.reset_value(1),.q(P02F0));
DFF_save_fm DFF_P48(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0300));
DFF_save_fm DFF_P49(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0310));
DFF_save_fm DFF_P50(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0320));
DFF_save_fm DFF_P51(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0330));
DFF_save_fm DFF_P52(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0340));
DFF_save_fm DFF_P53(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0350));
DFF_save_fm DFF_P54(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0360));
DFF_save_fm DFF_P55(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0370));
DFF_save_fm DFF_P56(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0380));
DFF_save_fm DFF_P57(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0390));
DFF_save_fm DFF_P58(.clk(clk),.rstn(rstn),.reset_value(1),.q(P03A0));
DFF_save_fm DFF_P59(.clk(clk),.rstn(rstn),.reset_value(0),.q(P03B0));
DFF_save_fm DFF_P60(.clk(clk),.rstn(rstn),.reset_value(0),.q(P03C0));
DFF_save_fm DFF_P61(.clk(clk),.rstn(rstn),.reset_value(1),.q(P03D0));
DFF_save_fm DFF_P62(.clk(clk),.rstn(rstn),.reset_value(1),.q(P03E0));
DFF_save_fm DFF_P63(.clk(clk),.rstn(rstn),.reset_value(1),.q(P03F0));
DFF_save_fm DFF_P64(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0400));
DFF_save_fm DFF_P65(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0410));
DFF_save_fm DFF_P66(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0420));
DFF_save_fm DFF_P67(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0430));
DFF_save_fm DFF_P68(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0440));
DFF_save_fm DFF_P69(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0450));
DFF_save_fm DFF_P70(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0460));
DFF_save_fm DFF_P71(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0470));
DFF_save_fm DFF_P72(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0480));
DFF_save_fm DFF_P73(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0490));
DFF_save_fm DFF_P74(.clk(clk),.rstn(rstn),.reset_value(1),.q(P04A0));
DFF_save_fm DFF_P75(.clk(clk),.rstn(rstn),.reset_value(1),.q(P04B0));
DFF_save_fm DFF_P76(.clk(clk),.rstn(rstn),.reset_value(0),.q(P04C0));
DFF_save_fm DFF_P77(.clk(clk),.rstn(rstn),.reset_value(1),.q(P04D0));
DFF_save_fm DFF_P78(.clk(clk),.rstn(rstn),.reset_value(1),.q(P04E0));
DFF_save_fm DFF_P79(.clk(clk),.rstn(rstn),.reset_value(1),.q(P04F0));
DFF_save_fm DFF_P80(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0500));
DFF_save_fm DFF_P81(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0510));
DFF_save_fm DFF_P82(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0520));
DFF_save_fm DFF_P83(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0530));
DFF_save_fm DFF_P84(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0540));
DFF_save_fm DFF_P85(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0550));
DFF_save_fm DFF_P86(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0560));
DFF_save_fm DFF_P87(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0570));
DFF_save_fm DFF_P88(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0580));
DFF_save_fm DFF_P89(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0590));
DFF_save_fm DFF_P90(.clk(clk),.rstn(rstn),.reset_value(1),.q(P05A0));
DFF_save_fm DFF_P91(.clk(clk),.rstn(rstn),.reset_value(1),.q(P05B0));
DFF_save_fm DFF_P92(.clk(clk),.rstn(rstn),.reset_value(1),.q(P05C0));
DFF_save_fm DFF_P93(.clk(clk),.rstn(rstn),.reset_value(1),.q(P05D0));
DFF_save_fm DFF_P94(.clk(clk),.rstn(rstn),.reset_value(1),.q(P05E0));
DFF_save_fm DFF_P95(.clk(clk),.rstn(rstn),.reset_value(1),.q(P05F0));
DFF_save_fm DFF_P96(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0600));
DFF_save_fm DFF_P97(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0610));
DFF_save_fm DFF_P98(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0620));
DFF_save_fm DFF_P99(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0630));
DFF_save_fm DFF_P100(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0640));
DFF_save_fm DFF_P101(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0650));
DFF_save_fm DFF_P102(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0660));
DFF_save_fm DFF_P103(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0670));
DFF_save_fm DFF_P104(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0680));
DFF_save_fm DFF_P105(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0690));
DFF_save_fm DFF_P106(.clk(clk),.rstn(rstn),.reset_value(1),.q(P06A0));
DFF_save_fm DFF_P107(.clk(clk),.rstn(rstn),.reset_value(1),.q(P06B0));
DFF_save_fm DFF_P108(.clk(clk),.rstn(rstn),.reset_value(1),.q(P06C0));
DFF_save_fm DFF_P109(.clk(clk),.rstn(rstn),.reset_value(1),.q(P06D0));
DFF_save_fm DFF_P110(.clk(clk),.rstn(rstn),.reset_value(1),.q(P06E0));
DFF_save_fm DFF_P111(.clk(clk),.rstn(rstn),.reset_value(1),.q(P06F0));
DFF_save_fm DFF_P112(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0700));
DFF_save_fm DFF_P113(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0710));
DFF_save_fm DFF_P114(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0720));
DFF_save_fm DFF_P115(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0730));
DFF_save_fm DFF_P116(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0740));
DFF_save_fm DFF_P117(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0750));
DFF_save_fm DFF_P118(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0760));
DFF_save_fm DFF_P119(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0770));
DFF_save_fm DFF_P120(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0780));
DFF_save_fm DFF_P121(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0790));
DFF_save_fm DFF_P122(.clk(clk),.rstn(rstn),.reset_value(1),.q(P07A0));
DFF_save_fm DFF_P123(.clk(clk),.rstn(rstn),.reset_value(1),.q(P07B0));
DFF_save_fm DFF_P124(.clk(clk),.rstn(rstn),.reset_value(1),.q(P07C0));
DFF_save_fm DFF_P125(.clk(clk),.rstn(rstn),.reset_value(1),.q(P07D0));
DFF_save_fm DFF_P126(.clk(clk),.rstn(rstn),.reset_value(1),.q(P07E0));
DFF_save_fm DFF_P127(.clk(clk),.rstn(rstn),.reset_value(1),.q(P07F0));
DFF_save_fm DFF_P128(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0800));
DFF_save_fm DFF_P129(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0810));
DFF_save_fm DFF_P130(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0820));
DFF_save_fm DFF_P131(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0830));
DFF_save_fm DFF_P132(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0840));
DFF_save_fm DFF_P133(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0850));
DFF_save_fm DFF_P134(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0860));
DFF_save_fm DFF_P135(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0870));
DFF_save_fm DFF_P136(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0880));
DFF_save_fm DFF_P137(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0890));
DFF_save_fm DFF_P138(.clk(clk),.rstn(rstn),.reset_value(1),.q(P08A0));
DFF_save_fm DFF_P139(.clk(clk),.rstn(rstn),.reset_value(1),.q(P08B0));
DFF_save_fm DFF_P140(.clk(clk),.rstn(rstn),.reset_value(1),.q(P08C0));
DFF_save_fm DFF_P141(.clk(clk),.rstn(rstn),.reset_value(1),.q(P08D0));
DFF_save_fm DFF_P142(.clk(clk),.rstn(rstn),.reset_value(1),.q(P08E0));
DFF_save_fm DFF_P143(.clk(clk),.rstn(rstn),.reset_value(1),.q(P08F0));
DFF_save_fm DFF_P144(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0900));
DFF_save_fm DFF_P145(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0910));
DFF_save_fm DFF_P146(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0920));
DFF_save_fm DFF_P147(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0930));
DFF_save_fm DFF_P148(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0940));
DFF_save_fm DFF_P149(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0950));
DFF_save_fm DFF_P150(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0960));
DFF_save_fm DFF_P151(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0970));
DFF_save_fm DFF_P152(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0980));
DFF_save_fm DFF_P153(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0990));
DFF_save_fm DFF_P154(.clk(clk),.rstn(rstn),.reset_value(1),.q(P09A0));
DFF_save_fm DFF_P155(.clk(clk),.rstn(rstn),.reset_value(1),.q(P09B0));
DFF_save_fm DFF_P156(.clk(clk),.rstn(rstn),.reset_value(1),.q(P09C0));
DFF_save_fm DFF_P157(.clk(clk),.rstn(rstn),.reset_value(1),.q(P09D0));
DFF_save_fm DFF_P158(.clk(clk),.rstn(rstn),.reset_value(1),.q(P09E0));
DFF_save_fm DFF_P159(.clk(clk),.rstn(rstn),.reset_value(1),.q(P09F0));
DFF_save_fm DFF_P160(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A00));
DFF_save_fm DFF_P161(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A10));
DFF_save_fm DFF_P162(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A20));
DFF_save_fm DFF_P163(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A30));
DFF_save_fm DFF_P164(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A40));
DFF_save_fm DFF_P165(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A50));
DFF_save_fm DFF_P166(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A60));
DFF_save_fm DFF_P167(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A70));
DFF_save_fm DFF_P168(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A80));
DFF_save_fm DFF_P169(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A90));
DFF_save_fm DFF_P170(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0AA0));
DFF_save_fm DFF_P171(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0AB0));
DFF_save_fm DFF_P172(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0AC0));
DFF_save_fm DFF_P173(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0AD0));
DFF_save_fm DFF_P174(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0AE0));
DFF_save_fm DFF_P175(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0AF0));
DFF_save_fm DFF_P176(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B00));
DFF_save_fm DFF_P177(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B10));
DFF_save_fm DFF_P178(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B20));
DFF_save_fm DFF_P179(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B30));
DFF_save_fm DFF_P180(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B40));
DFF_save_fm DFF_P181(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B50));
DFF_save_fm DFF_P182(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B60));
DFF_save_fm DFF_P183(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B70));
DFF_save_fm DFF_P184(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B80));
DFF_save_fm DFF_P185(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B90));
DFF_save_fm DFF_P186(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0BA0));
DFF_save_fm DFF_P187(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0BB0));
DFF_save_fm DFF_P188(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0BC0));
DFF_save_fm DFF_P189(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0BD0));
DFF_save_fm DFF_P190(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0BE0));
DFF_save_fm DFF_P191(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0BF0));
DFF_save_fm DFF_P192(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C00));
DFF_save_fm DFF_P193(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C10));
DFF_save_fm DFF_P194(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C20));
DFF_save_fm DFF_P195(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C30));
DFF_save_fm DFF_P196(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C40));
DFF_save_fm DFF_P197(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C50));
DFF_save_fm DFF_P198(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C60));
DFF_save_fm DFF_P199(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C70));
DFF_save_fm DFF_P200(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C80));
DFF_save_fm DFF_P201(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C90));
DFF_save_fm DFF_P202(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0CA0));
DFF_save_fm DFF_P203(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0CB0));
DFF_save_fm DFF_P204(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0CC0));
DFF_save_fm DFF_P205(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0CD0));
DFF_save_fm DFF_P206(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0CE0));
DFF_save_fm DFF_P207(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0CF0));
DFF_save_fm DFF_P208(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D00));
DFF_save_fm DFF_P209(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D10));
DFF_save_fm DFF_P210(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D20));
DFF_save_fm DFF_P211(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D30));
DFF_save_fm DFF_P212(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D40));
DFF_save_fm DFF_P213(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D50));
DFF_save_fm DFF_P214(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D60));
DFF_save_fm DFF_P215(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D70));
DFF_save_fm DFF_P216(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D80));
DFF_save_fm DFF_P217(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D90));
DFF_save_fm DFF_P218(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0DA0));
DFF_save_fm DFF_P219(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0DB0));
DFF_save_fm DFF_P220(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0DC0));
DFF_save_fm DFF_P221(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0DD0));
DFF_save_fm DFF_P222(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0DE0));
DFF_save_fm DFF_P223(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0DF0));
DFF_save_fm DFF_P224(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E00));
DFF_save_fm DFF_P225(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E10));
DFF_save_fm DFF_P226(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E20));
DFF_save_fm DFF_P227(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E30));
DFF_save_fm DFF_P228(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E40));
DFF_save_fm DFF_P229(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E50));
DFF_save_fm DFF_P230(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E60));
DFF_save_fm DFF_P231(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E70));
DFF_save_fm DFF_P232(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E80));
DFF_save_fm DFF_P233(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E90));
DFF_save_fm DFF_P234(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0EA0));
DFF_save_fm DFF_P235(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0EB0));
DFF_save_fm DFF_P236(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0EC0));
DFF_save_fm DFF_P237(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0ED0));
DFF_save_fm DFF_P238(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0EE0));
DFF_save_fm DFF_P239(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0EF0));
DFF_save_fm DFF_P240(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F00));
DFF_save_fm DFF_P241(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F10));
DFF_save_fm DFF_P242(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F20));
DFF_save_fm DFF_P243(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F30));
DFF_save_fm DFF_P244(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F40));
DFF_save_fm DFF_P245(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F50));
DFF_save_fm DFF_P246(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F60));
DFF_save_fm DFF_P247(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F70));
DFF_save_fm DFF_P248(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F80));
DFF_save_fm DFF_P249(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F90));
DFF_save_fm DFF_P250(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0FA0));
DFF_save_fm DFF_P251(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0FB0));
DFF_save_fm DFF_P252(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0FC0));
DFF_save_fm DFF_P253(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0FD0));
DFF_save_fm DFF_P254(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0FE0));
DFF_save_fm DFF_P255(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0FF0));
DFF_save_fm DFF_P256(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0001));
DFF_save_fm DFF_P257(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0011));
DFF_save_fm DFF_P258(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0021));
DFF_save_fm DFF_P259(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0031));
DFF_save_fm DFF_P260(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0041));
DFF_save_fm DFF_P261(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0051));
DFF_save_fm DFF_P262(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0061));
DFF_save_fm DFF_P263(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0071));
DFF_save_fm DFF_P264(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0081));
DFF_save_fm DFF_P265(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0091));
DFF_save_fm DFF_P266(.clk(clk),.rstn(rstn),.reset_value(1),.q(P00A1));
DFF_save_fm DFF_P267(.clk(clk),.rstn(rstn),.reset_value(1),.q(P00B1));
DFF_save_fm DFF_P268(.clk(clk),.rstn(rstn),.reset_value(1),.q(P00C1));
DFF_save_fm DFF_P269(.clk(clk),.rstn(rstn),.reset_value(1),.q(P00D1));
DFF_save_fm DFF_P270(.clk(clk),.rstn(rstn),.reset_value(1),.q(P00E1));
DFF_save_fm DFF_P271(.clk(clk),.rstn(rstn),.reset_value(1),.q(P00F1));
DFF_save_fm DFF_P272(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0101));
DFF_save_fm DFF_P273(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0111));
DFF_save_fm DFF_P274(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0121));
DFF_save_fm DFF_P275(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0131));
DFF_save_fm DFF_P276(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0141));
DFF_save_fm DFF_P277(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0151));
DFF_save_fm DFF_P278(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0161));
DFF_save_fm DFF_P279(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0171));
DFF_save_fm DFF_P280(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0181));
DFF_save_fm DFF_P281(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0191));
DFF_save_fm DFF_P282(.clk(clk),.rstn(rstn),.reset_value(0),.q(P01A1));
DFF_save_fm DFF_P283(.clk(clk),.rstn(rstn),.reset_value(0),.q(P01B1));
DFF_save_fm DFF_P284(.clk(clk),.rstn(rstn),.reset_value(0),.q(P01C1));
DFF_save_fm DFF_P285(.clk(clk),.rstn(rstn),.reset_value(1),.q(P01D1));
DFF_save_fm DFF_P286(.clk(clk),.rstn(rstn),.reset_value(1),.q(P01E1));
DFF_save_fm DFF_P287(.clk(clk),.rstn(rstn),.reset_value(1),.q(P01F1));
DFF_save_fm DFF_P288(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0201));
DFF_save_fm DFF_P289(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0211));
DFF_save_fm DFF_P290(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0221));
DFF_save_fm DFF_P291(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0231));
DFF_save_fm DFF_P292(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0241));
DFF_save_fm DFF_P293(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0251));
DFF_save_fm DFF_P294(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0261));
DFF_save_fm DFF_P295(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0271));
DFF_save_fm DFF_P296(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0281));
DFF_save_fm DFF_P297(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0291));
DFF_save_fm DFF_P298(.clk(clk),.rstn(rstn),.reset_value(0),.q(P02A1));
DFF_save_fm DFF_P299(.clk(clk),.rstn(rstn),.reset_value(0),.q(P02B1));
DFF_save_fm DFF_P300(.clk(clk),.rstn(rstn),.reset_value(0),.q(P02C1));
DFF_save_fm DFF_P301(.clk(clk),.rstn(rstn),.reset_value(1),.q(P02D1));
DFF_save_fm DFF_P302(.clk(clk),.rstn(rstn),.reset_value(1),.q(P02E1));
DFF_save_fm DFF_P303(.clk(clk),.rstn(rstn),.reset_value(1),.q(P02F1));
DFF_save_fm DFF_P304(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0301));
DFF_save_fm DFF_P305(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0311));
DFF_save_fm DFF_P306(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0321));
DFF_save_fm DFF_P307(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0331));
DFF_save_fm DFF_P308(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0341));
DFF_save_fm DFF_P309(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0351));
DFF_save_fm DFF_P310(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0361));
DFF_save_fm DFF_P311(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0371));
DFF_save_fm DFF_P312(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0381));
DFF_save_fm DFF_P313(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0391));
DFF_save_fm DFF_P314(.clk(clk),.rstn(rstn),.reset_value(0),.q(P03A1));
DFF_save_fm DFF_P315(.clk(clk),.rstn(rstn),.reset_value(0),.q(P03B1));
DFF_save_fm DFF_P316(.clk(clk),.rstn(rstn),.reset_value(0),.q(P03C1));
DFF_save_fm DFF_P317(.clk(clk),.rstn(rstn),.reset_value(1),.q(P03D1));
DFF_save_fm DFF_P318(.clk(clk),.rstn(rstn),.reset_value(1),.q(P03E1));
DFF_save_fm DFF_P319(.clk(clk),.rstn(rstn),.reset_value(1),.q(P03F1));
DFF_save_fm DFF_P320(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0401));
DFF_save_fm DFF_P321(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0411));
DFF_save_fm DFF_P322(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0421));
DFF_save_fm DFF_P323(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0431));
DFF_save_fm DFF_P324(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0441));
DFF_save_fm DFF_P325(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0451));
DFF_save_fm DFF_P326(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0461));
DFF_save_fm DFF_P327(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0471));
DFF_save_fm DFF_P328(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0481));
DFF_save_fm DFF_P329(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0491));
DFF_save_fm DFF_P330(.clk(clk),.rstn(rstn),.reset_value(0),.q(P04A1));
DFF_save_fm DFF_P331(.clk(clk),.rstn(rstn),.reset_value(0),.q(P04B1));
DFF_save_fm DFF_P332(.clk(clk),.rstn(rstn),.reset_value(0),.q(P04C1));
DFF_save_fm DFF_P333(.clk(clk),.rstn(rstn),.reset_value(1),.q(P04D1));
DFF_save_fm DFF_P334(.clk(clk),.rstn(rstn),.reset_value(1),.q(P04E1));
DFF_save_fm DFF_P335(.clk(clk),.rstn(rstn),.reset_value(1),.q(P04F1));
DFF_save_fm DFF_P336(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0501));
DFF_save_fm DFF_P337(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0511));
DFF_save_fm DFF_P338(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0521));
DFF_save_fm DFF_P339(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0531));
DFF_save_fm DFF_P340(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0541));
DFF_save_fm DFF_P341(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0551));
DFF_save_fm DFF_P342(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0561));
DFF_save_fm DFF_P343(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0571));
DFF_save_fm DFF_P344(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0581));
DFF_save_fm DFF_P345(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0591));
DFF_save_fm DFF_P346(.clk(clk),.rstn(rstn),.reset_value(1),.q(P05A1));
DFF_save_fm DFF_P347(.clk(clk),.rstn(rstn),.reset_value(0),.q(P05B1));
DFF_save_fm DFF_P348(.clk(clk),.rstn(rstn),.reset_value(0),.q(P05C1));
DFF_save_fm DFF_P349(.clk(clk),.rstn(rstn),.reset_value(1),.q(P05D1));
DFF_save_fm DFF_P350(.clk(clk),.rstn(rstn),.reset_value(1),.q(P05E1));
DFF_save_fm DFF_P351(.clk(clk),.rstn(rstn),.reset_value(1),.q(P05F1));
DFF_save_fm DFF_P352(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0601));
DFF_save_fm DFF_P353(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0611));
DFF_save_fm DFF_P354(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0621));
DFF_save_fm DFF_P355(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0631));
DFF_save_fm DFF_P356(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0641));
DFF_save_fm DFF_P357(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0651));
DFF_save_fm DFF_P358(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0661));
DFF_save_fm DFF_P359(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0671));
DFF_save_fm DFF_P360(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0681));
DFF_save_fm DFF_P361(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0691));
DFF_save_fm DFF_P362(.clk(clk),.rstn(rstn),.reset_value(1),.q(P06A1));
DFF_save_fm DFF_P363(.clk(clk),.rstn(rstn),.reset_value(1),.q(P06B1));
DFF_save_fm DFF_P364(.clk(clk),.rstn(rstn),.reset_value(1),.q(P06C1));
DFF_save_fm DFF_P365(.clk(clk),.rstn(rstn),.reset_value(1),.q(P06D1));
DFF_save_fm DFF_P366(.clk(clk),.rstn(rstn),.reset_value(1),.q(P06E1));
DFF_save_fm DFF_P367(.clk(clk),.rstn(rstn),.reset_value(1),.q(P06F1));
DFF_save_fm DFF_P368(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0701));
DFF_save_fm DFF_P369(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0711));
DFF_save_fm DFF_P370(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0721));
DFF_save_fm DFF_P371(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0731));
DFF_save_fm DFF_P372(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0741));
DFF_save_fm DFF_P373(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0751));
DFF_save_fm DFF_P374(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0761));
DFF_save_fm DFF_P375(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0771));
DFF_save_fm DFF_P376(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0781));
DFF_save_fm DFF_P377(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0791));
DFF_save_fm DFF_P378(.clk(clk),.rstn(rstn),.reset_value(1),.q(P07A1));
DFF_save_fm DFF_P379(.clk(clk),.rstn(rstn),.reset_value(1),.q(P07B1));
DFF_save_fm DFF_P380(.clk(clk),.rstn(rstn),.reset_value(1),.q(P07C1));
DFF_save_fm DFF_P381(.clk(clk),.rstn(rstn),.reset_value(1),.q(P07D1));
DFF_save_fm DFF_P382(.clk(clk),.rstn(rstn),.reset_value(1),.q(P07E1));
DFF_save_fm DFF_P383(.clk(clk),.rstn(rstn),.reset_value(1),.q(P07F1));
DFF_save_fm DFF_P384(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0801));
DFF_save_fm DFF_P385(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0811));
DFF_save_fm DFF_P386(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0821));
DFF_save_fm DFF_P387(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0831));
DFF_save_fm DFF_P388(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0841));
DFF_save_fm DFF_P389(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0851));
DFF_save_fm DFF_P390(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0861));
DFF_save_fm DFF_P391(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0871));
DFF_save_fm DFF_P392(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0881));
DFF_save_fm DFF_P393(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0891));
DFF_save_fm DFF_P394(.clk(clk),.rstn(rstn),.reset_value(1),.q(P08A1));
DFF_save_fm DFF_P395(.clk(clk),.rstn(rstn),.reset_value(1),.q(P08B1));
DFF_save_fm DFF_P396(.clk(clk),.rstn(rstn),.reset_value(1),.q(P08C1));
DFF_save_fm DFF_P397(.clk(clk),.rstn(rstn),.reset_value(1),.q(P08D1));
DFF_save_fm DFF_P398(.clk(clk),.rstn(rstn),.reset_value(1),.q(P08E1));
DFF_save_fm DFF_P399(.clk(clk),.rstn(rstn),.reset_value(1),.q(P08F1));
DFF_save_fm DFF_P400(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0901));
DFF_save_fm DFF_P401(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0911));
DFF_save_fm DFF_P402(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0921));
DFF_save_fm DFF_P403(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0931));
DFF_save_fm DFF_P404(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0941));
DFF_save_fm DFF_P405(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0951));
DFF_save_fm DFF_P406(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0961));
DFF_save_fm DFF_P407(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0971));
DFF_save_fm DFF_P408(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0981));
DFF_save_fm DFF_P409(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0991));
DFF_save_fm DFF_P410(.clk(clk),.rstn(rstn),.reset_value(1),.q(P09A1));
DFF_save_fm DFF_P411(.clk(clk),.rstn(rstn),.reset_value(1),.q(P09B1));
DFF_save_fm DFF_P412(.clk(clk),.rstn(rstn),.reset_value(1),.q(P09C1));
DFF_save_fm DFF_P413(.clk(clk),.rstn(rstn),.reset_value(1),.q(P09D1));
DFF_save_fm DFF_P414(.clk(clk),.rstn(rstn),.reset_value(1),.q(P09E1));
DFF_save_fm DFF_P415(.clk(clk),.rstn(rstn),.reset_value(1),.q(P09F1));
DFF_save_fm DFF_P416(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A01));
DFF_save_fm DFF_P417(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A11));
DFF_save_fm DFF_P418(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A21));
DFF_save_fm DFF_P419(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A31));
DFF_save_fm DFF_P420(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A41));
DFF_save_fm DFF_P421(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A51));
DFF_save_fm DFF_P422(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A61));
DFF_save_fm DFF_P423(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A71));
DFF_save_fm DFF_P424(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A81));
DFF_save_fm DFF_P425(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A91));
DFF_save_fm DFF_P426(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0AA1));
DFF_save_fm DFF_P427(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0AB1));
DFF_save_fm DFF_P428(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0AC1));
DFF_save_fm DFF_P429(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0AD1));
DFF_save_fm DFF_P430(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0AE1));
DFF_save_fm DFF_P431(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0AF1));
DFF_save_fm DFF_P432(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B01));
DFF_save_fm DFF_P433(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B11));
DFF_save_fm DFF_P434(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B21));
DFF_save_fm DFF_P435(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B31));
DFF_save_fm DFF_P436(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B41));
DFF_save_fm DFF_P437(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B51));
DFF_save_fm DFF_P438(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B61));
DFF_save_fm DFF_P439(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B71));
DFF_save_fm DFF_P440(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B81));
DFF_save_fm DFF_P441(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B91));
DFF_save_fm DFF_P442(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0BA1));
DFF_save_fm DFF_P443(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0BB1));
DFF_save_fm DFF_P444(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0BC1));
DFF_save_fm DFF_P445(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0BD1));
DFF_save_fm DFF_P446(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0BE1));
DFF_save_fm DFF_P447(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0BF1));
DFF_save_fm DFF_P448(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C01));
DFF_save_fm DFF_P449(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C11));
DFF_save_fm DFF_P450(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C21));
DFF_save_fm DFF_P451(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C31));
DFF_save_fm DFF_P452(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C41));
DFF_save_fm DFF_P453(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C51));
DFF_save_fm DFF_P454(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C61));
DFF_save_fm DFF_P455(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C71));
DFF_save_fm DFF_P456(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C81));
DFF_save_fm DFF_P457(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C91));
DFF_save_fm DFF_P458(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0CA1));
DFF_save_fm DFF_P459(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0CB1));
DFF_save_fm DFF_P460(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0CC1));
DFF_save_fm DFF_P461(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0CD1));
DFF_save_fm DFF_P462(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0CE1));
DFF_save_fm DFF_P463(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0CF1));
DFF_save_fm DFF_P464(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D01));
DFF_save_fm DFF_P465(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D11));
DFF_save_fm DFF_P466(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D21));
DFF_save_fm DFF_P467(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D31));
DFF_save_fm DFF_P468(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D41));
DFF_save_fm DFF_P469(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0D51));
DFF_save_fm DFF_P470(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D61));
DFF_save_fm DFF_P471(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D71));
DFF_save_fm DFF_P472(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D81));
DFF_save_fm DFF_P473(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D91));
DFF_save_fm DFF_P474(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0DA1));
DFF_save_fm DFF_P475(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0DB1));
DFF_save_fm DFF_P476(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0DC1));
DFF_save_fm DFF_P477(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0DD1));
DFF_save_fm DFF_P478(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0DE1));
DFF_save_fm DFF_P479(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0DF1));
DFF_save_fm DFF_P480(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E01));
DFF_save_fm DFF_P481(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E11));
DFF_save_fm DFF_P482(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E21));
DFF_save_fm DFF_P483(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E31));
DFF_save_fm DFF_P484(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E41));
DFF_save_fm DFF_P485(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0E51));
DFF_save_fm DFF_P486(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0E61));
DFF_save_fm DFF_P487(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E71));
DFF_save_fm DFF_P488(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E81));
DFF_save_fm DFF_P489(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0E91));
DFF_save_fm DFF_P490(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0EA1));
DFF_save_fm DFF_P491(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0EB1));
DFF_save_fm DFF_P492(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0EC1));
DFF_save_fm DFF_P493(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0ED1));
DFF_save_fm DFF_P494(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0EE1));
DFF_save_fm DFF_P495(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0EF1));
DFF_save_fm DFF_P496(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F01));
DFF_save_fm DFF_P497(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F11));
DFF_save_fm DFF_P498(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F21));
DFF_save_fm DFF_P499(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F31));
DFF_save_fm DFF_P500(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F41));
DFF_save_fm DFF_P501(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F51));
DFF_save_fm DFF_P502(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F61));
DFF_save_fm DFF_P503(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F71));
DFF_save_fm DFF_P504(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F81));
DFF_save_fm DFF_P505(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F91));
DFF_save_fm DFF_P506(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0FA1));
DFF_save_fm DFF_P507(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0FB1));
DFF_save_fm DFF_P508(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0FC1));
DFF_save_fm DFF_P509(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0FD1));
DFF_save_fm DFF_P510(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0FE1));
DFF_save_fm DFF_P511(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0FF1));
DFF_save_fm DFF_P512(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0002));
DFF_save_fm DFF_P513(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0012));
DFF_save_fm DFF_P514(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0022));
DFF_save_fm DFF_P515(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0032));
DFF_save_fm DFF_P516(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0042));
DFF_save_fm DFF_P517(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0052));
DFF_save_fm DFF_P518(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0062));
DFF_save_fm DFF_P519(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0072));
DFF_save_fm DFF_P520(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0082));
DFF_save_fm DFF_P521(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0092));
DFF_save_fm DFF_P522(.clk(clk),.rstn(rstn),.reset_value(1),.q(P00A2));
DFF_save_fm DFF_P523(.clk(clk),.rstn(rstn),.reset_value(1),.q(P00B2));
DFF_save_fm DFF_P524(.clk(clk),.rstn(rstn),.reset_value(1),.q(P00C2));
DFF_save_fm DFF_P525(.clk(clk),.rstn(rstn),.reset_value(1),.q(P00D2));
DFF_save_fm DFF_P526(.clk(clk),.rstn(rstn),.reset_value(1),.q(P00E2));
DFF_save_fm DFF_P527(.clk(clk),.rstn(rstn),.reset_value(1),.q(P00F2));
DFF_save_fm DFF_P528(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0102));
DFF_save_fm DFF_P529(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0112));
DFF_save_fm DFF_P530(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0122));
DFF_save_fm DFF_P531(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0132));
DFF_save_fm DFF_P532(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0142));
DFF_save_fm DFF_P533(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0152));
DFF_save_fm DFF_P534(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0162));
DFF_save_fm DFF_P535(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0172));
DFF_save_fm DFF_P536(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0182));
DFF_save_fm DFF_P537(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0192));
DFF_save_fm DFF_P538(.clk(clk),.rstn(rstn),.reset_value(0),.q(P01A2));
DFF_save_fm DFF_P539(.clk(clk),.rstn(rstn),.reset_value(0),.q(P01B2));
DFF_save_fm DFF_P540(.clk(clk),.rstn(rstn),.reset_value(0),.q(P01C2));
DFF_save_fm DFF_P541(.clk(clk),.rstn(rstn),.reset_value(1),.q(P01D2));
DFF_save_fm DFF_P542(.clk(clk),.rstn(rstn),.reset_value(1),.q(P01E2));
DFF_save_fm DFF_P543(.clk(clk),.rstn(rstn),.reset_value(1),.q(P01F2));
DFF_save_fm DFF_P544(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0202));
DFF_save_fm DFF_P545(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0212));
DFF_save_fm DFF_P546(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0222));
DFF_save_fm DFF_P547(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0232));
DFF_save_fm DFF_P548(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0242));
DFF_save_fm DFF_P549(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0252));
DFF_save_fm DFF_P550(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0262));
DFF_save_fm DFF_P551(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0272));
DFF_save_fm DFF_P552(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0282));
DFF_save_fm DFF_P553(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0292));
DFF_save_fm DFF_P554(.clk(clk),.rstn(rstn),.reset_value(0),.q(P02A2));
DFF_save_fm DFF_P555(.clk(clk),.rstn(rstn),.reset_value(0),.q(P02B2));
DFF_save_fm DFF_P556(.clk(clk),.rstn(rstn),.reset_value(0),.q(P02C2));
DFF_save_fm DFF_P557(.clk(clk),.rstn(rstn),.reset_value(1),.q(P02D2));
DFF_save_fm DFF_P558(.clk(clk),.rstn(rstn),.reset_value(1),.q(P02E2));
DFF_save_fm DFF_P559(.clk(clk),.rstn(rstn),.reset_value(1),.q(P02F2));
DFF_save_fm DFF_P560(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0302));
DFF_save_fm DFF_P561(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0312));
DFF_save_fm DFF_P562(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0322));
DFF_save_fm DFF_P563(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0332));
DFF_save_fm DFF_P564(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0342));
DFF_save_fm DFF_P565(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0352));
DFF_save_fm DFF_P566(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0362));
DFF_save_fm DFF_P567(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0372));
DFF_save_fm DFF_P568(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0382));
DFF_save_fm DFF_P569(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0392));
DFF_save_fm DFF_P570(.clk(clk),.rstn(rstn),.reset_value(0),.q(P03A2));
DFF_save_fm DFF_P571(.clk(clk),.rstn(rstn),.reset_value(0),.q(P03B2));
DFF_save_fm DFF_P572(.clk(clk),.rstn(rstn),.reset_value(0),.q(P03C2));
DFF_save_fm DFF_P573(.clk(clk),.rstn(rstn),.reset_value(1),.q(P03D2));
DFF_save_fm DFF_P574(.clk(clk),.rstn(rstn),.reset_value(1),.q(P03E2));
DFF_save_fm DFF_P575(.clk(clk),.rstn(rstn),.reset_value(1),.q(P03F2));
DFF_save_fm DFF_P576(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0402));
DFF_save_fm DFF_P577(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0412));
DFF_save_fm DFF_P578(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0422));
DFF_save_fm DFF_P579(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0432));
DFF_save_fm DFF_P580(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0442));
DFF_save_fm DFF_P581(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0452));
DFF_save_fm DFF_P582(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0462));
DFF_save_fm DFF_P583(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0472));
DFF_save_fm DFF_P584(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0482));
DFF_save_fm DFF_P585(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0492));
DFF_save_fm DFF_P586(.clk(clk),.rstn(rstn),.reset_value(0),.q(P04A2));
DFF_save_fm DFF_P587(.clk(clk),.rstn(rstn),.reset_value(0),.q(P04B2));
DFF_save_fm DFF_P588(.clk(clk),.rstn(rstn),.reset_value(0),.q(P04C2));
DFF_save_fm DFF_P589(.clk(clk),.rstn(rstn),.reset_value(1),.q(P04D2));
DFF_save_fm DFF_P590(.clk(clk),.rstn(rstn),.reset_value(1),.q(P04E2));
DFF_save_fm DFF_P591(.clk(clk),.rstn(rstn),.reset_value(1),.q(P04F2));
DFF_save_fm DFF_P592(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0502));
DFF_save_fm DFF_P593(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0512));
DFF_save_fm DFF_P594(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0522));
DFF_save_fm DFF_P595(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0532));
DFF_save_fm DFF_P596(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0542));
DFF_save_fm DFF_P597(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0552));
DFF_save_fm DFF_P598(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0562));
DFF_save_fm DFF_P599(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0572));
DFF_save_fm DFF_P600(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0582));
DFF_save_fm DFF_P601(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0592));
DFF_save_fm DFF_P602(.clk(clk),.rstn(rstn),.reset_value(0),.q(P05A2));
DFF_save_fm DFF_P603(.clk(clk),.rstn(rstn),.reset_value(0),.q(P05B2));
DFF_save_fm DFF_P604(.clk(clk),.rstn(rstn),.reset_value(0),.q(P05C2));
DFF_save_fm DFF_P605(.clk(clk),.rstn(rstn),.reset_value(1),.q(P05D2));
DFF_save_fm DFF_P606(.clk(clk),.rstn(rstn),.reset_value(1),.q(P05E2));
DFF_save_fm DFF_P607(.clk(clk),.rstn(rstn),.reset_value(1),.q(P05F2));
DFF_save_fm DFF_P608(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0602));
DFF_save_fm DFF_P609(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0612));
DFF_save_fm DFF_P610(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0622));
DFF_save_fm DFF_P611(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0632));
DFF_save_fm DFF_P612(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0642));
DFF_save_fm DFF_P613(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0652));
DFF_save_fm DFF_P614(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0662));
DFF_save_fm DFF_P615(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0672));
DFF_save_fm DFF_P616(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0682));
DFF_save_fm DFF_P617(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0692));
DFF_save_fm DFF_P618(.clk(clk),.rstn(rstn),.reset_value(1),.q(P06A2));
DFF_save_fm DFF_P619(.clk(clk),.rstn(rstn),.reset_value(0),.q(P06B2));
DFF_save_fm DFF_P620(.clk(clk),.rstn(rstn),.reset_value(0),.q(P06C2));
DFF_save_fm DFF_P621(.clk(clk),.rstn(rstn),.reset_value(1),.q(P06D2));
DFF_save_fm DFF_P622(.clk(clk),.rstn(rstn),.reset_value(1),.q(P06E2));
DFF_save_fm DFF_P623(.clk(clk),.rstn(rstn),.reset_value(1),.q(P06F2));
DFF_save_fm DFF_P624(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0702));
DFF_save_fm DFF_P625(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0712));
DFF_save_fm DFF_P626(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0722));
DFF_save_fm DFF_P627(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0732));
DFF_save_fm DFF_P628(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0742));
DFF_save_fm DFF_P629(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0752));
DFF_save_fm DFF_P630(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0762));
DFF_save_fm DFF_P631(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0772));
DFF_save_fm DFF_P632(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0782));
DFF_save_fm DFF_P633(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0792));
DFF_save_fm DFF_P634(.clk(clk),.rstn(rstn),.reset_value(1),.q(P07A2));
DFF_save_fm DFF_P635(.clk(clk),.rstn(rstn),.reset_value(1),.q(P07B2));
DFF_save_fm DFF_P636(.clk(clk),.rstn(rstn),.reset_value(0),.q(P07C2));
DFF_save_fm DFF_P637(.clk(clk),.rstn(rstn),.reset_value(1),.q(P07D2));
DFF_save_fm DFF_P638(.clk(clk),.rstn(rstn),.reset_value(1),.q(P07E2));
DFF_save_fm DFF_P639(.clk(clk),.rstn(rstn),.reset_value(1),.q(P07F2));
DFF_save_fm DFF_P640(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0802));
DFF_save_fm DFF_P641(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0812));
DFF_save_fm DFF_P642(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0822));
DFF_save_fm DFF_P643(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0832));
DFF_save_fm DFF_P644(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0842));
DFF_save_fm DFF_P645(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0852));
DFF_save_fm DFF_P646(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0862));
DFF_save_fm DFF_P647(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0872));
DFF_save_fm DFF_P648(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0882));
DFF_save_fm DFF_P649(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0892));
DFF_save_fm DFF_P650(.clk(clk),.rstn(rstn),.reset_value(1),.q(P08A2));
DFF_save_fm DFF_P651(.clk(clk),.rstn(rstn),.reset_value(1),.q(P08B2));
DFF_save_fm DFF_P652(.clk(clk),.rstn(rstn),.reset_value(1),.q(P08C2));
DFF_save_fm DFF_P653(.clk(clk),.rstn(rstn),.reset_value(1),.q(P08D2));
DFF_save_fm DFF_P654(.clk(clk),.rstn(rstn),.reset_value(1),.q(P08E2));
DFF_save_fm DFF_P655(.clk(clk),.rstn(rstn),.reset_value(1),.q(P08F2));
DFF_save_fm DFF_P656(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0902));
DFF_save_fm DFF_P657(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0912));
DFF_save_fm DFF_P658(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0922));
DFF_save_fm DFF_P659(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0932));
DFF_save_fm DFF_P660(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0942));
DFF_save_fm DFF_P661(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0952));
DFF_save_fm DFF_P662(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0962));
DFF_save_fm DFF_P663(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0972));
DFF_save_fm DFF_P664(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0982));
DFF_save_fm DFF_P665(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0992));
DFF_save_fm DFF_P666(.clk(clk),.rstn(rstn),.reset_value(1),.q(P09A2));
DFF_save_fm DFF_P667(.clk(clk),.rstn(rstn),.reset_value(1),.q(P09B2));
DFF_save_fm DFF_P668(.clk(clk),.rstn(rstn),.reset_value(1),.q(P09C2));
DFF_save_fm DFF_P669(.clk(clk),.rstn(rstn),.reset_value(1),.q(P09D2));
DFF_save_fm DFF_P670(.clk(clk),.rstn(rstn),.reset_value(1),.q(P09E2));
DFF_save_fm DFF_P671(.clk(clk),.rstn(rstn),.reset_value(1),.q(P09F2));
DFF_save_fm DFF_P672(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A02));
DFF_save_fm DFF_P673(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A12));
DFF_save_fm DFF_P674(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A22));
DFF_save_fm DFF_P675(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A32));
DFF_save_fm DFF_P676(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A42));
DFF_save_fm DFF_P677(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A52));
DFF_save_fm DFF_P678(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A62));
DFF_save_fm DFF_P679(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A72));
DFF_save_fm DFF_P680(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A82));
DFF_save_fm DFF_P681(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0A92));
DFF_save_fm DFF_P682(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0AA2));
DFF_save_fm DFF_P683(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0AB2));
DFF_save_fm DFF_P684(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0AC2));
DFF_save_fm DFF_P685(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0AD2));
DFF_save_fm DFF_P686(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0AE2));
DFF_save_fm DFF_P687(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0AF2));
DFF_save_fm DFF_P688(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B02));
DFF_save_fm DFF_P689(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B12));
DFF_save_fm DFF_P690(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B22));
DFF_save_fm DFF_P691(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B32));
DFF_save_fm DFF_P692(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B42));
DFF_save_fm DFF_P693(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B52));
DFF_save_fm DFF_P694(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B62));
DFF_save_fm DFF_P695(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B72));
DFF_save_fm DFF_P696(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B82));
DFF_save_fm DFF_P697(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0B92));
DFF_save_fm DFF_P698(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0BA2));
DFF_save_fm DFF_P699(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0BB2));
DFF_save_fm DFF_P700(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0BC2));
DFF_save_fm DFF_P701(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0BD2));
DFF_save_fm DFF_P702(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0BE2));
DFF_save_fm DFF_P703(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0BF2));
DFF_save_fm DFF_P704(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C02));
DFF_save_fm DFF_P705(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C12));
DFF_save_fm DFF_P706(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C22));
DFF_save_fm DFF_P707(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C32));
DFF_save_fm DFF_P708(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C42));
DFF_save_fm DFF_P709(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C52));
DFF_save_fm DFF_P710(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C62));
DFF_save_fm DFF_P711(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C72));
DFF_save_fm DFF_P712(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C82));
DFF_save_fm DFF_P713(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0C92));
DFF_save_fm DFF_P714(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0CA2));
DFF_save_fm DFF_P715(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0CB2));
DFF_save_fm DFF_P716(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0CC2));
DFF_save_fm DFF_P717(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0CD2));
DFF_save_fm DFF_P718(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0CE2));
DFF_save_fm DFF_P719(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0CF2));
DFF_save_fm DFF_P720(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D02));
DFF_save_fm DFF_P721(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D12));
DFF_save_fm DFF_P722(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D22));
DFF_save_fm DFF_P723(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D32));
DFF_save_fm DFF_P724(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D42));
DFF_save_fm DFF_P725(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0D52));
DFF_save_fm DFF_P726(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0D62));
DFF_save_fm DFF_P727(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D72));
DFF_save_fm DFF_P728(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0D82));
DFF_save_fm DFF_P729(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0D92));
DFF_save_fm DFF_P730(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0DA2));
DFF_save_fm DFF_P731(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0DB2));
DFF_save_fm DFF_P732(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0DC2));
DFF_save_fm DFF_P733(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0DD2));
DFF_save_fm DFF_P734(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0DE2));
DFF_save_fm DFF_P735(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0DF2));
DFF_save_fm DFF_P736(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E02));
DFF_save_fm DFF_P737(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E12));
DFF_save_fm DFF_P738(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E22));
DFF_save_fm DFF_P739(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E32));
DFF_save_fm DFF_P740(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0E42));
DFF_save_fm DFF_P741(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0E52));
DFF_save_fm DFF_P742(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0E62));
DFF_save_fm DFF_P743(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0E72));
DFF_save_fm DFF_P744(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0E82));
DFF_save_fm DFF_P745(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0E92));
DFF_save_fm DFF_P746(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0EA2));
DFF_save_fm DFF_P747(.clk(clk),.rstn(rstn),.reset_value(0),.q(P0EB2));
DFF_save_fm DFF_P748(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0EC2));
DFF_save_fm DFF_P749(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0ED2));
DFF_save_fm DFF_P750(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0EE2));
DFF_save_fm DFF_P751(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0EF2));
DFF_save_fm DFF_P752(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F02));
DFF_save_fm DFF_P753(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F12));
DFF_save_fm DFF_P754(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F22));
DFF_save_fm DFF_P755(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F32));
DFF_save_fm DFF_P756(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F42));
DFF_save_fm DFF_P757(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F52));
DFF_save_fm DFF_P758(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F62));
DFF_save_fm DFF_P759(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F72));
DFF_save_fm DFF_P760(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F82));
DFF_save_fm DFF_P761(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0F92));
DFF_save_fm DFF_P762(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0FA2));
DFF_save_fm DFF_P763(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0FB2));
DFF_save_fm DFF_P764(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0FC2));
DFF_save_fm DFF_P765(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0FD2));
DFF_save_fm DFF_P766(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0FE2));
DFF_save_fm DFF_P767(.clk(clk),.rstn(rstn),.reset_value(1),.q(P0FF2));
DFF_save_fm DFF_W0(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00000));
DFF_save_fm DFF_W1(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00010));
DFF_save_fm DFF_W2(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00020));
DFF_save_fm DFF_W3(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00100));
DFF_save_fm DFF_W4(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00110));
DFF_save_fm DFF_W5(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00120));
DFF_save_fm DFF_W6(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00200));
DFF_save_fm DFF_W7(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00210));
DFF_save_fm DFF_W8(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00220));
DFF_save_fm DFF_W9(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00001));
DFF_save_fm DFF_W10(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00011));
DFF_save_fm DFF_W11(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00021));
DFF_save_fm DFF_W12(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00101));
DFF_save_fm DFF_W13(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00111));
DFF_save_fm DFF_W14(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00121));
DFF_save_fm DFF_W15(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00201));
DFF_save_fm DFF_W16(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00211));
DFF_save_fm DFF_W17(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00221));
DFF_save_fm DFF_W18(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00002));
DFF_save_fm DFF_W19(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00012));
DFF_save_fm DFF_W20(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00022));
DFF_save_fm DFF_W21(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00102));
DFF_save_fm DFF_W22(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00112));
DFF_save_fm DFF_W23(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00122));
DFF_save_fm DFF_W24(.clk(clk),.rstn(rstn),.reset_value(0),.q(W00202));
DFF_save_fm DFF_W25(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00212));
DFF_save_fm DFF_W26(.clk(clk),.rstn(rstn),.reset_value(1),.q(W00222));
DFF_save_fm DFF_W27(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01000));
DFF_save_fm DFF_W28(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01010));
DFF_save_fm DFF_W29(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01020));
DFF_save_fm DFF_W30(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01100));
DFF_save_fm DFF_W31(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01110));
DFF_save_fm DFF_W32(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01120));
DFF_save_fm DFF_W33(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01200));
DFF_save_fm DFF_W34(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01210));
DFF_save_fm DFF_W35(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01220));
DFF_save_fm DFF_W36(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01001));
DFF_save_fm DFF_W37(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01011));
DFF_save_fm DFF_W38(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01021));
DFF_save_fm DFF_W39(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01101));
DFF_save_fm DFF_W40(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01111));
DFF_save_fm DFF_W41(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01121));
DFF_save_fm DFF_W42(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01201));
DFF_save_fm DFF_W43(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01211));
DFF_save_fm DFF_W44(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01221));
DFF_save_fm DFF_W45(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01002));
DFF_save_fm DFF_W46(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01012));
DFF_save_fm DFF_W47(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01022));
DFF_save_fm DFF_W48(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01102));
DFF_save_fm DFF_W49(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01112));
DFF_save_fm DFF_W50(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01122));
DFF_save_fm DFF_W51(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01202));
DFF_save_fm DFF_W52(.clk(clk),.rstn(rstn),.reset_value(1),.q(W01212));
DFF_save_fm DFF_W53(.clk(clk),.rstn(rstn),.reset_value(0),.q(W01222));
DFF_save_fm DFF_W54(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02000));
DFF_save_fm DFF_W55(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02010));
DFF_save_fm DFF_W56(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02020));
DFF_save_fm DFF_W57(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02100));
DFF_save_fm DFF_W58(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02110));
DFF_save_fm DFF_W59(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02120));
DFF_save_fm DFF_W60(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02200));
DFF_save_fm DFF_W61(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02210));
DFF_save_fm DFF_W62(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02220));
DFF_save_fm DFF_W63(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02001));
DFF_save_fm DFF_W64(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02011));
DFF_save_fm DFF_W65(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02021));
DFF_save_fm DFF_W66(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02101));
DFF_save_fm DFF_W67(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02111));
DFF_save_fm DFF_W68(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02121));
DFF_save_fm DFF_W69(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02201));
DFF_save_fm DFF_W70(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02211));
DFF_save_fm DFF_W71(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02221));
DFF_save_fm DFF_W72(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02002));
DFF_save_fm DFF_W73(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02012));
DFF_save_fm DFF_W74(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02022));
DFF_save_fm DFF_W75(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02102));
DFF_save_fm DFF_W76(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02112));
DFF_save_fm DFF_W77(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02122));
DFF_save_fm DFF_W78(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02202));
DFF_save_fm DFF_W79(.clk(clk),.rstn(rstn),.reset_value(1),.q(W02212));
DFF_save_fm DFF_W80(.clk(clk),.rstn(rstn),.reset_value(0),.q(W02222));
ninexnine_unit ninexnine_unit_0(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00000)
);

ninexnine_unit ninexnine_unit_1(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01000)
);

ninexnine_unit ninexnine_unit_2(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02000)
);

assign C0000=c00000+c01000+c02000;
assign A0000=(C0000>=0)?1:0;

ninexnine_unit ninexnine_unit_3(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00010)
);

ninexnine_unit ninexnine_unit_4(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01010)
);

ninexnine_unit ninexnine_unit_5(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02010)
);

assign C0010=c00010+c01010+c02010;
assign A0010=(C0010>=0)?1:0;

ninexnine_unit ninexnine_unit_6(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00020)
);

ninexnine_unit ninexnine_unit_7(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01020)
);

ninexnine_unit ninexnine_unit_8(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02020)
);

assign C0020=c00020+c01020+c02020;
assign A0020=(C0020>=0)?1:0;

ninexnine_unit ninexnine_unit_9(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00030)
);

ninexnine_unit ninexnine_unit_10(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01030)
);

ninexnine_unit ninexnine_unit_11(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02030)
);

assign C0030=c00030+c01030+c02030;
assign A0030=(C0030>=0)?1:0;

ninexnine_unit ninexnine_unit_12(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00040)
);

ninexnine_unit ninexnine_unit_13(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01040)
);

ninexnine_unit ninexnine_unit_14(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02040)
);

assign C0040=c00040+c01040+c02040;
assign A0040=(C0040>=0)?1:0;

ninexnine_unit ninexnine_unit_15(
				.clk(clk),
				.rstn(rstn),
				.a0(P0050),
				.a1(P0060),
				.a2(P0070),
				.a3(P0150),
				.a4(P0160),
				.a5(P0170),
				.a6(P0250),
				.a7(P0260),
				.a8(P0270),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00050)
);

ninexnine_unit ninexnine_unit_16(
				.clk(clk),
				.rstn(rstn),
				.a0(P0051),
				.a1(P0061),
				.a2(P0071),
				.a3(P0151),
				.a4(P0161),
				.a5(P0171),
				.a6(P0251),
				.a7(P0261),
				.a8(P0271),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01050)
);

ninexnine_unit ninexnine_unit_17(
				.clk(clk),
				.rstn(rstn),
				.a0(P0052),
				.a1(P0062),
				.a2(P0072),
				.a3(P0152),
				.a4(P0162),
				.a5(P0172),
				.a6(P0252),
				.a7(P0262),
				.a8(P0272),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02050)
);

assign C0050=c00050+c01050+c02050;
assign A0050=(C0050>=0)?1:0;

ninexnine_unit ninexnine_unit_18(
				.clk(clk),
				.rstn(rstn),
				.a0(P0060),
				.a1(P0070),
				.a2(P0080),
				.a3(P0160),
				.a4(P0170),
				.a5(P0180),
				.a6(P0260),
				.a7(P0270),
				.a8(P0280),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00060)
);

ninexnine_unit ninexnine_unit_19(
				.clk(clk),
				.rstn(rstn),
				.a0(P0061),
				.a1(P0071),
				.a2(P0081),
				.a3(P0161),
				.a4(P0171),
				.a5(P0181),
				.a6(P0261),
				.a7(P0271),
				.a8(P0281),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01060)
);

ninexnine_unit ninexnine_unit_20(
				.clk(clk),
				.rstn(rstn),
				.a0(P0062),
				.a1(P0072),
				.a2(P0082),
				.a3(P0162),
				.a4(P0172),
				.a5(P0182),
				.a6(P0262),
				.a7(P0272),
				.a8(P0282),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02060)
);

assign C0060=c00060+c01060+c02060;
assign A0060=(C0060>=0)?1:0;

ninexnine_unit ninexnine_unit_21(
				.clk(clk),
				.rstn(rstn),
				.a0(P0070),
				.a1(P0080),
				.a2(P0090),
				.a3(P0170),
				.a4(P0180),
				.a5(P0190),
				.a6(P0270),
				.a7(P0280),
				.a8(P0290),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00070)
);

ninexnine_unit ninexnine_unit_22(
				.clk(clk),
				.rstn(rstn),
				.a0(P0071),
				.a1(P0081),
				.a2(P0091),
				.a3(P0171),
				.a4(P0181),
				.a5(P0191),
				.a6(P0271),
				.a7(P0281),
				.a8(P0291),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01070)
);

ninexnine_unit ninexnine_unit_23(
				.clk(clk),
				.rstn(rstn),
				.a0(P0072),
				.a1(P0082),
				.a2(P0092),
				.a3(P0172),
				.a4(P0182),
				.a5(P0192),
				.a6(P0272),
				.a7(P0282),
				.a8(P0292),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02070)
);

assign C0070=c00070+c01070+c02070;
assign A0070=(C0070>=0)?1:0;

ninexnine_unit ninexnine_unit_24(
				.clk(clk),
				.rstn(rstn),
				.a0(P0080),
				.a1(P0090),
				.a2(P00A0),
				.a3(P0180),
				.a4(P0190),
				.a5(P01A0),
				.a6(P0280),
				.a7(P0290),
				.a8(P02A0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00080)
);

ninexnine_unit ninexnine_unit_25(
				.clk(clk),
				.rstn(rstn),
				.a0(P0081),
				.a1(P0091),
				.a2(P00A1),
				.a3(P0181),
				.a4(P0191),
				.a5(P01A1),
				.a6(P0281),
				.a7(P0291),
				.a8(P02A1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01080)
);

ninexnine_unit ninexnine_unit_26(
				.clk(clk),
				.rstn(rstn),
				.a0(P0082),
				.a1(P0092),
				.a2(P00A2),
				.a3(P0182),
				.a4(P0192),
				.a5(P01A2),
				.a6(P0282),
				.a7(P0292),
				.a8(P02A2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02080)
);

assign C0080=c00080+c01080+c02080;
assign A0080=(C0080>=0)?1:0;

ninexnine_unit ninexnine_unit_27(
				.clk(clk),
				.rstn(rstn),
				.a0(P0090),
				.a1(P00A0),
				.a2(P00B0),
				.a3(P0190),
				.a4(P01A0),
				.a5(P01B0),
				.a6(P0290),
				.a7(P02A0),
				.a8(P02B0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00090)
);

ninexnine_unit ninexnine_unit_28(
				.clk(clk),
				.rstn(rstn),
				.a0(P0091),
				.a1(P00A1),
				.a2(P00B1),
				.a3(P0191),
				.a4(P01A1),
				.a5(P01B1),
				.a6(P0291),
				.a7(P02A1),
				.a8(P02B1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01090)
);

ninexnine_unit ninexnine_unit_29(
				.clk(clk),
				.rstn(rstn),
				.a0(P0092),
				.a1(P00A2),
				.a2(P00B2),
				.a3(P0192),
				.a4(P01A2),
				.a5(P01B2),
				.a6(P0292),
				.a7(P02A2),
				.a8(P02B2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02090)
);

assign C0090=c00090+c01090+c02090;
assign A0090=(C0090>=0)?1:0;

ninexnine_unit ninexnine_unit_30(
				.clk(clk),
				.rstn(rstn),
				.a0(P00A0),
				.a1(P00B0),
				.a2(P00C0),
				.a3(P01A0),
				.a4(P01B0),
				.a5(P01C0),
				.a6(P02A0),
				.a7(P02B0),
				.a8(P02C0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c000A0)
);

ninexnine_unit ninexnine_unit_31(
				.clk(clk),
				.rstn(rstn),
				.a0(P00A1),
				.a1(P00B1),
				.a2(P00C1),
				.a3(P01A1),
				.a4(P01B1),
				.a5(P01C1),
				.a6(P02A1),
				.a7(P02B1),
				.a8(P02C1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c010A0)
);

ninexnine_unit ninexnine_unit_32(
				.clk(clk),
				.rstn(rstn),
				.a0(P00A2),
				.a1(P00B2),
				.a2(P00C2),
				.a3(P01A2),
				.a4(P01B2),
				.a5(P01C2),
				.a6(P02A2),
				.a7(P02B2),
				.a8(P02C2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c020A0)
);

assign C00A0=c000A0+c010A0+c020A0;
assign A00A0=(C00A0>=0)?1:0;

ninexnine_unit ninexnine_unit_33(
				.clk(clk),
				.rstn(rstn),
				.a0(P00B0),
				.a1(P00C0),
				.a2(P00D0),
				.a3(P01B0),
				.a4(P01C0),
				.a5(P01D0),
				.a6(P02B0),
				.a7(P02C0),
				.a8(P02D0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c000B0)
);

ninexnine_unit ninexnine_unit_34(
				.clk(clk),
				.rstn(rstn),
				.a0(P00B1),
				.a1(P00C1),
				.a2(P00D1),
				.a3(P01B1),
				.a4(P01C1),
				.a5(P01D1),
				.a6(P02B1),
				.a7(P02C1),
				.a8(P02D1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c010B0)
);

ninexnine_unit ninexnine_unit_35(
				.clk(clk),
				.rstn(rstn),
				.a0(P00B2),
				.a1(P00C2),
				.a2(P00D2),
				.a3(P01B2),
				.a4(P01C2),
				.a5(P01D2),
				.a6(P02B2),
				.a7(P02C2),
				.a8(P02D2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c020B0)
);

assign C00B0=c000B0+c010B0+c020B0;
assign A00B0=(C00B0>=0)?1:0;

ninexnine_unit ninexnine_unit_36(
				.clk(clk),
				.rstn(rstn),
				.a0(P00C0),
				.a1(P00D0),
				.a2(P00E0),
				.a3(P01C0),
				.a4(P01D0),
				.a5(P01E0),
				.a6(P02C0),
				.a7(P02D0),
				.a8(P02E0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c000C0)
);

ninexnine_unit ninexnine_unit_37(
				.clk(clk),
				.rstn(rstn),
				.a0(P00C1),
				.a1(P00D1),
				.a2(P00E1),
				.a3(P01C1),
				.a4(P01D1),
				.a5(P01E1),
				.a6(P02C1),
				.a7(P02D1),
				.a8(P02E1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c010C0)
);

ninexnine_unit ninexnine_unit_38(
				.clk(clk),
				.rstn(rstn),
				.a0(P00C2),
				.a1(P00D2),
				.a2(P00E2),
				.a3(P01C2),
				.a4(P01D2),
				.a5(P01E2),
				.a6(P02C2),
				.a7(P02D2),
				.a8(P02E2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c020C0)
);

assign C00C0=c000C0+c010C0+c020C0;
assign A00C0=(C00C0>=0)?1:0;

ninexnine_unit ninexnine_unit_39(
				.clk(clk),
				.rstn(rstn),
				.a0(P00D0),
				.a1(P00E0),
				.a2(P00F0),
				.a3(P01D0),
				.a4(P01E0),
				.a5(P01F0),
				.a6(P02D0),
				.a7(P02E0),
				.a8(P02F0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c000D0)
);

ninexnine_unit ninexnine_unit_40(
				.clk(clk),
				.rstn(rstn),
				.a0(P00D1),
				.a1(P00E1),
				.a2(P00F1),
				.a3(P01D1),
				.a4(P01E1),
				.a5(P01F1),
				.a6(P02D1),
				.a7(P02E1),
				.a8(P02F1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c010D0)
);

ninexnine_unit ninexnine_unit_41(
				.clk(clk),
				.rstn(rstn),
				.a0(P00D2),
				.a1(P00E2),
				.a2(P00F2),
				.a3(P01D2),
				.a4(P01E2),
				.a5(P01F2),
				.a6(P02D2),
				.a7(P02E2),
				.a8(P02F2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c020D0)
);

assign C00D0=c000D0+c010D0+c020D0;
assign A00D0=(C00D0>=0)?1:0;

ninexnine_unit ninexnine_unit_42(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00100)
);

ninexnine_unit ninexnine_unit_43(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01100)
);

ninexnine_unit ninexnine_unit_44(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02100)
);

assign C0100=c00100+c01100+c02100;
assign A0100=(C0100>=0)?1:0;

ninexnine_unit ninexnine_unit_45(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00110)
);

ninexnine_unit ninexnine_unit_46(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01110)
);

ninexnine_unit ninexnine_unit_47(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02110)
);

assign C0110=c00110+c01110+c02110;
assign A0110=(C0110>=0)?1:0;

ninexnine_unit ninexnine_unit_48(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00120)
);

ninexnine_unit ninexnine_unit_49(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01120)
);

ninexnine_unit ninexnine_unit_50(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02120)
);

assign C0120=c00120+c01120+c02120;
assign A0120=(C0120>=0)?1:0;

ninexnine_unit ninexnine_unit_51(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00130)
);

ninexnine_unit ninexnine_unit_52(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01130)
);

ninexnine_unit ninexnine_unit_53(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02130)
);

assign C0130=c00130+c01130+c02130;
assign A0130=(C0130>=0)?1:0;

ninexnine_unit ninexnine_unit_54(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00140)
);

ninexnine_unit ninexnine_unit_55(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01140)
);

ninexnine_unit ninexnine_unit_56(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02140)
);

assign C0140=c00140+c01140+c02140;
assign A0140=(C0140>=0)?1:0;

ninexnine_unit ninexnine_unit_57(
				.clk(clk),
				.rstn(rstn),
				.a0(P0150),
				.a1(P0160),
				.a2(P0170),
				.a3(P0250),
				.a4(P0260),
				.a5(P0270),
				.a6(P0350),
				.a7(P0360),
				.a8(P0370),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00150)
);

ninexnine_unit ninexnine_unit_58(
				.clk(clk),
				.rstn(rstn),
				.a0(P0151),
				.a1(P0161),
				.a2(P0171),
				.a3(P0251),
				.a4(P0261),
				.a5(P0271),
				.a6(P0351),
				.a7(P0361),
				.a8(P0371),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01150)
);

ninexnine_unit ninexnine_unit_59(
				.clk(clk),
				.rstn(rstn),
				.a0(P0152),
				.a1(P0162),
				.a2(P0172),
				.a3(P0252),
				.a4(P0262),
				.a5(P0272),
				.a6(P0352),
				.a7(P0362),
				.a8(P0372),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02150)
);

assign C0150=c00150+c01150+c02150;
assign A0150=(C0150>=0)?1:0;

ninexnine_unit ninexnine_unit_60(
				.clk(clk),
				.rstn(rstn),
				.a0(P0160),
				.a1(P0170),
				.a2(P0180),
				.a3(P0260),
				.a4(P0270),
				.a5(P0280),
				.a6(P0360),
				.a7(P0370),
				.a8(P0380),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00160)
);

ninexnine_unit ninexnine_unit_61(
				.clk(clk),
				.rstn(rstn),
				.a0(P0161),
				.a1(P0171),
				.a2(P0181),
				.a3(P0261),
				.a4(P0271),
				.a5(P0281),
				.a6(P0361),
				.a7(P0371),
				.a8(P0381),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01160)
);

ninexnine_unit ninexnine_unit_62(
				.clk(clk),
				.rstn(rstn),
				.a0(P0162),
				.a1(P0172),
				.a2(P0182),
				.a3(P0262),
				.a4(P0272),
				.a5(P0282),
				.a6(P0362),
				.a7(P0372),
				.a8(P0382),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02160)
);

assign C0160=c00160+c01160+c02160;
assign A0160=(C0160>=0)?1:0;

ninexnine_unit ninexnine_unit_63(
				.clk(clk),
				.rstn(rstn),
				.a0(P0170),
				.a1(P0180),
				.a2(P0190),
				.a3(P0270),
				.a4(P0280),
				.a5(P0290),
				.a6(P0370),
				.a7(P0380),
				.a8(P0390),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00170)
);

ninexnine_unit ninexnine_unit_64(
				.clk(clk),
				.rstn(rstn),
				.a0(P0171),
				.a1(P0181),
				.a2(P0191),
				.a3(P0271),
				.a4(P0281),
				.a5(P0291),
				.a6(P0371),
				.a7(P0381),
				.a8(P0391),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01170)
);

ninexnine_unit ninexnine_unit_65(
				.clk(clk),
				.rstn(rstn),
				.a0(P0172),
				.a1(P0182),
				.a2(P0192),
				.a3(P0272),
				.a4(P0282),
				.a5(P0292),
				.a6(P0372),
				.a7(P0382),
				.a8(P0392),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02170)
);

assign C0170=c00170+c01170+c02170;
assign A0170=(C0170>=0)?1:0;

ninexnine_unit ninexnine_unit_66(
				.clk(clk),
				.rstn(rstn),
				.a0(P0180),
				.a1(P0190),
				.a2(P01A0),
				.a3(P0280),
				.a4(P0290),
				.a5(P02A0),
				.a6(P0380),
				.a7(P0390),
				.a8(P03A0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00180)
);

ninexnine_unit ninexnine_unit_67(
				.clk(clk),
				.rstn(rstn),
				.a0(P0181),
				.a1(P0191),
				.a2(P01A1),
				.a3(P0281),
				.a4(P0291),
				.a5(P02A1),
				.a6(P0381),
				.a7(P0391),
				.a8(P03A1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01180)
);

ninexnine_unit ninexnine_unit_68(
				.clk(clk),
				.rstn(rstn),
				.a0(P0182),
				.a1(P0192),
				.a2(P01A2),
				.a3(P0282),
				.a4(P0292),
				.a5(P02A2),
				.a6(P0382),
				.a7(P0392),
				.a8(P03A2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02180)
);

assign C0180=c00180+c01180+c02180;
assign A0180=(C0180>=0)?1:0;

ninexnine_unit ninexnine_unit_69(
				.clk(clk),
				.rstn(rstn),
				.a0(P0190),
				.a1(P01A0),
				.a2(P01B0),
				.a3(P0290),
				.a4(P02A0),
				.a5(P02B0),
				.a6(P0390),
				.a7(P03A0),
				.a8(P03B0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00190)
);

ninexnine_unit ninexnine_unit_70(
				.clk(clk),
				.rstn(rstn),
				.a0(P0191),
				.a1(P01A1),
				.a2(P01B1),
				.a3(P0291),
				.a4(P02A1),
				.a5(P02B1),
				.a6(P0391),
				.a7(P03A1),
				.a8(P03B1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01190)
);

ninexnine_unit ninexnine_unit_71(
				.clk(clk),
				.rstn(rstn),
				.a0(P0192),
				.a1(P01A2),
				.a2(P01B2),
				.a3(P0292),
				.a4(P02A2),
				.a5(P02B2),
				.a6(P0392),
				.a7(P03A2),
				.a8(P03B2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02190)
);

assign C0190=c00190+c01190+c02190;
assign A0190=(C0190>=0)?1:0;

ninexnine_unit ninexnine_unit_72(
				.clk(clk),
				.rstn(rstn),
				.a0(P01A0),
				.a1(P01B0),
				.a2(P01C0),
				.a3(P02A0),
				.a4(P02B0),
				.a5(P02C0),
				.a6(P03A0),
				.a7(P03B0),
				.a8(P03C0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c001A0)
);

ninexnine_unit ninexnine_unit_73(
				.clk(clk),
				.rstn(rstn),
				.a0(P01A1),
				.a1(P01B1),
				.a2(P01C1),
				.a3(P02A1),
				.a4(P02B1),
				.a5(P02C1),
				.a6(P03A1),
				.a7(P03B1),
				.a8(P03C1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c011A0)
);

ninexnine_unit ninexnine_unit_74(
				.clk(clk),
				.rstn(rstn),
				.a0(P01A2),
				.a1(P01B2),
				.a2(P01C2),
				.a3(P02A2),
				.a4(P02B2),
				.a5(P02C2),
				.a6(P03A2),
				.a7(P03B2),
				.a8(P03C2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c021A0)
);

assign C01A0=c001A0+c011A0+c021A0;
assign A01A0=(C01A0>=0)?1:0;

ninexnine_unit ninexnine_unit_75(
				.clk(clk),
				.rstn(rstn),
				.a0(P01B0),
				.a1(P01C0),
				.a2(P01D0),
				.a3(P02B0),
				.a4(P02C0),
				.a5(P02D0),
				.a6(P03B0),
				.a7(P03C0),
				.a8(P03D0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c001B0)
);

ninexnine_unit ninexnine_unit_76(
				.clk(clk),
				.rstn(rstn),
				.a0(P01B1),
				.a1(P01C1),
				.a2(P01D1),
				.a3(P02B1),
				.a4(P02C1),
				.a5(P02D1),
				.a6(P03B1),
				.a7(P03C1),
				.a8(P03D1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c011B0)
);

ninexnine_unit ninexnine_unit_77(
				.clk(clk),
				.rstn(rstn),
				.a0(P01B2),
				.a1(P01C2),
				.a2(P01D2),
				.a3(P02B2),
				.a4(P02C2),
				.a5(P02D2),
				.a6(P03B2),
				.a7(P03C2),
				.a8(P03D2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c021B0)
);

assign C01B0=c001B0+c011B0+c021B0;
assign A01B0=(C01B0>=0)?1:0;

ninexnine_unit ninexnine_unit_78(
				.clk(clk),
				.rstn(rstn),
				.a0(P01C0),
				.a1(P01D0),
				.a2(P01E0),
				.a3(P02C0),
				.a4(P02D0),
				.a5(P02E0),
				.a6(P03C0),
				.a7(P03D0),
				.a8(P03E0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c001C0)
);

ninexnine_unit ninexnine_unit_79(
				.clk(clk),
				.rstn(rstn),
				.a0(P01C1),
				.a1(P01D1),
				.a2(P01E1),
				.a3(P02C1),
				.a4(P02D1),
				.a5(P02E1),
				.a6(P03C1),
				.a7(P03D1),
				.a8(P03E1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c011C0)
);

ninexnine_unit ninexnine_unit_80(
				.clk(clk),
				.rstn(rstn),
				.a0(P01C2),
				.a1(P01D2),
				.a2(P01E2),
				.a3(P02C2),
				.a4(P02D2),
				.a5(P02E2),
				.a6(P03C2),
				.a7(P03D2),
				.a8(P03E2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c021C0)
);

assign C01C0=c001C0+c011C0+c021C0;
assign A01C0=(C01C0>=0)?1:0;

ninexnine_unit ninexnine_unit_81(
				.clk(clk),
				.rstn(rstn),
				.a0(P01D0),
				.a1(P01E0),
				.a2(P01F0),
				.a3(P02D0),
				.a4(P02E0),
				.a5(P02F0),
				.a6(P03D0),
				.a7(P03E0),
				.a8(P03F0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c001D0)
);

ninexnine_unit ninexnine_unit_82(
				.clk(clk),
				.rstn(rstn),
				.a0(P01D1),
				.a1(P01E1),
				.a2(P01F1),
				.a3(P02D1),
				.a4(P02E1),
				.a5(P02F1),
				.a6(P03D1),
				.a7(P03E1),
				.a8(P03F1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c011D0)
);

ninexnine_unit ninexnine_unit_83(
				.clk(clk),
				.rstn(rstn),
				.a0(P01D2),
				.a1(P01E2),
				.a2(P01F2),
				.a3(P02D2),
				.a4(P02E2),
				.a5(P02F2),
				.a6(P03D2),
				.a7(P03E2),
				.a8(P03F2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c021D0)
);

assign C01D0=c001D0+c011D0+c021D0;
assign A01D0=(C01D0>=0)?1:0;

ninexnine_unit ninexnine_unit_84(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00200)
);

ninexnine_unit ninexnine_unit_85(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01200)
);

ninexnine_unit ninexnine_unit_86(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02200)
);

assign C0200=c00200+c01200+c02200;
assign A0200=(C0200>=0)?1:0;

ninexnine_unit ninexnine_unit_87(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00210)
);

ninexnine_unit ninexnine_unit_88(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01210)
);

ninexnine_unit ninexnine_unit_89(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02210)
);

assign C0210=c00210+c01210+c02210;
assign A0210=(C0210>=0)?1:0;

ninexnine_unit ninexnine_unit_90(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00220)
);

ninexnine_unit ninexnine_unit_91(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01220)
);

ninexnine_unit ninexnine_unit_92(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02220)
);

assign C0220=c00220+c01220+c02220;
assign A0220=(C0220>=0)?1:0;

ninexnine_unit ninexnine_unit_93(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00230)
);

ninexnine_unit ninexnine_unit_94(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01230)
);

ninexnine_unit ninexnine_unit_95(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02230)
);

assign C0230=c00230+c01230+c02230;
assign A0230=(C0230>=0)?1:0;

ninexnine_unit ninexnine_unit_96(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00240)
);

ninexnine_unit ninexnine_unit_97(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01240)
);

ninexnine_unit ninexnine_unit_98(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02240)
);

assign C0240=c00240+c01240+c02240;
assign A0240=(C0240>=0)?1:0;

ninexnine_unit ninexnine_unit_99(
				.clk(clk),
				.rstn(rstn),
				.a0(P0250),
				.a1(P0260),
				.a2(P0270),
				.a3(P0350),
				.a4(P0360),
				.a5(P0370),
				.a6(P0450),
				.a7(P0460),
				.a8(P0470),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00250)
);

ninexnine_unit ninexnine_unit_100(
				.clk(clk),
				.rstn(rstn),
				.a0(P0251),
				.a1(P0261),
				.a2(P0271),
				.a3(P0351),
				.a4(P0361),
				.a5(P0371),
				.a6(P0451),
				.a7(P0461),
				.a8(P0471),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01250)
);

ninexnine_unit ninexnine_unit_101(
				.clk(clk),
				.rstn(rstn),
				.a0(P0252),
				.a1(P0262),
				.a2(P0272),
				.a3(P0352),
				.a4(P0362),
				.a5(P0372),
				.a6(P0452),
				.a7(P0462),
				.a8(P0472),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02250)
);

assign C0250=c00250+c01250+c02250;
assign A0250=(C0250>=0)?1:0;

ninexnine_unit ninexnine_unit_102(
				.clk(clk),
				.rstn(rstn),
				.a0(P0260),
				.a1(P0270),
				.a2(P0280),
				.a3(P0360),
				.a4(P0370),
				.a5(P0380),
				.a6(P0460),
				.a7(P0470),
				.a8(P0480),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00260)
);

ninexnine_unit ninexnine_unit_103(
				.clk(clk),
				.rstn(rstn),
				.a0(P0261),
				.a1(P0271),
				.a2(P0281),
				.a3(P0361),
				.a4(P0371),
				.a5(P0381),
				.a6(P0461),
				.a7(P0471),
				.a8(P0481),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01260)
);

ninexnine_unit ninexnine_unit_104(
				.clk(clk),
				.rstn(rstn),
				.a0(P0262),
				.a1(P0272),
				.a2(P0282),
				.a3(P0362),
				.a4(P0372),
				.a5(P0382),
				.a6(P0462),
				.a7(P0472),
				.a8(P0482),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02260)
);

assign C0260=c00260+c01260+c02260;
assign A0260=(C0260>=0)?1:0;

ninexnine_unit ninexnine_unit_105(
				.clk(clk),
				.rstn(rstn),
				.a0(P0270),
				.a1(P0280),
				.a2(P0290),
				.a3(P0370),
				.a4(P0380),
				.a5(P0390),
				.a6(P0470),
				.a7(P0480),
				.a8(P0490),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00270)
);

ninexnine_unit ninexnine_unit_106(
				.clk(clk),
				.rstn(rstn),
				.a0(P0271),
				.a1(P0281),
				.a2(P0291),
				.a3(P0371),
				.a4(P0381),
				.a5(P0391),
				.a6(P0471),
				.a7(P0481),
				.a8(P0491),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01270)
);

ninexnine_unit ninexnine_unit_107(
				.clk(clk),
				.rstn(rstn),
				.a0(P0272),
				.a1(P0282),
				.a2(P0292),
				.a3(P0372),
				.a4(P0382),
				.a5(P0392),
				.a6(P0472),
				.a7(P0482),
				.a8(P0492),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02270)
);

assign C0270=c00270+c01270+c02270;
assign A0270=(C0270>=0)?1:0;

ninexnine_unit ninexnine_unit_108(
				.clk(clk),
				.rstn(rstn),
				.a0(P0280),
				.a1(P0290),
				.a2(P02A0),
				.a3(P0380),
				.a4(P0390),
				.a5(P03A0),
				.a6(P0480),
				.a7(P0490),
				.a8(P04A0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00280)
);

ninexnine_unit ninexnine_unit_109(
				.clk(clk),
				.rstn(rstn),
				.a0(P0281),
				.a1(P0291),
				.a2(P02A1),
				.a3(P0381),
				.a4(P0391),
				.a5(P03A1),
				.a6(P0481),
				.a7(P0491),
				.a8(P04A1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01280)
);

ninexnine_unit ninexnine_unit_110(
				.clk(clk),
				.rstn(rstn),
				.a0(P0282),
				.a1(P0292),
				.a2(P02A2),
				.a3(P0382),
				.a4(P0392),
				.a5(P03A2),
				.a6(P0482),
				.a7(P0492),
				.a8(P04A2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02280)
);

assign C0280=c00280+c01280+c02280;
assign A0280=(C0280>=0)?1:0;

ninexnine_unit ninexnine_unit_111(
				.clk(clk),
				.rstn(rstn),
				.a0(P0290),
				.a1(P02A0),
				.a2(P02B0),
				.a3(P0390),
				.a4(P03A0),
				.a5(P03B0),
				.a6(P0490),
				.a7(P04A0),
				.a8(P04B0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00290)
);

ninexnine_unit ninexnine_unit_112(
				.clk(clk),
				.rstn(rstn),
				.a0(P0291),
				.a1(P02A1),
				.a2(P02B1),
				.a3(P0391),
				.a4(P03A1),
				.a5(P03B1),
				.a6(P0491),
				.a7(P04A1),
				.a8(P04B1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01290)
);

ninexnine_unit ninexnine_unit_113(
				.clk(clk),
				.rstn(rstn),
				.a0(P0292),
				.a1(P02A2),
				.a2(P02B2),
				.a3(P0392),
				.a4(P03A2),
				.a5(P03B2),
				.a6(P0492),
				.a7(P04A2),
				.a8(P04B2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02290)
);

assign C0290=c00290+c01290+c02290;
assign A0290=(C0290>=0)?1:0;

ninexnine_unit ninexnine_unit_114(
				.clk(clk),
				.rstn(rstn),
				.a0(P02A0),
				.a1(P02B0),
				.a2(P02C0),
				.a3(P03A0),
				.a4(P03B0),
				.a5(P03C0),
				.a6(P04A0),
				.a7(P04B0),
				.a8(P04C0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c002A0)
);

ninexnine_unit ninexnine_unit_115(
				.clk(clk),
				.rstn(rstn),
				.a0(P02A1),
				.a1(P02B1),
				.a2(P02C1),
				.a3(P03A1),
				.a4(P03B1),
				.a5(P03C1),
				.a6(P04A1),
				.a7(P04B1),
				.a8(P04C1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c012A0)
);

ninexnine_unit ninexnine_unit_116(
				.clk(clk),
				.rstn(rstn),
				.a0(P02A2),
				.a1(P02B2),
				.a2(P02C2),
				.a3(P03A2),
				.a4(P03B2),
				.a5(P03C2),
				.a6(P04A2),
				.a7(P04B2),
				.a8(P04C2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c022A0)
);

assign C02A0=c002A0+c012A0+c022A0;
assign A02A0=(C02A0>=0)?1:0;

ninexnine_unit ninexnine_unit_117(
				.clk(clk),
				.rstn(rstn),
				.a0(P02B0),
				.a1(P02C0),
				.a2(P02D0),
				.a3(P03B0),
				.a4(P03C0),
				.a5(P03D0),
				.a6(P04B0),
				.a7(P04C0),
				.a8(P04D0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c002B0)
);

ninexnine_unit ninexnine_unit_118(
				.clk(clk),
				.rstn(rstn),
				.a0(P02B1),
				.a1(P02C1),
				.a2(P02D1),
				.a3(P03B1),
				.a4(P03C1),
				.a5(P03D1),
				.a6(P04B1),
				.a7(P04C1),
				.a8(P04D1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c012B0)
);

ninexnine_unit ninexnine_unit_119(
				.clk(clk),
				.rstn(rstn),
				.a0(P02B2),
				.a1(P02C2),
				.a2(P02D2),
				.a3(P03B2),
				.a4(P03C2),
				.a5(P03D2),
				.a6(P04B2),
				.a7(P04C2),
				.a8(P04D2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c022B0)
);

assign C02B0=c002B0+c012B0+c022B0;
assign A02B0=(C02B0>=0)?1:0;

ninexnine_unit ninexnine_unit_120(
				.clk(clk),
				.rstn(rstn),
				.a0(P02C0),
				.a1(P02D0),
				.a2(P02E0),
				.a3(P03C0),
				.a4(P03D0),
				.a5(P03E0),
				.a6(P04C0),
				.a7(P04D0),
				.a8(P04E0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c002C0)
);

ninexnine_unit ninexnine_unit_121(
				.clk(clk),
				.rstn(rstn),
				.a0(P02C1),
				.a1(P02D1),
				.a2(P02E1),
				.a3(P03C1),
				.a4(P03D1),
				.a5(P03E1),
				.a6(P04C1),
				.a7(P04D1),
				.a8(P04E1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c012C0)
);

ninexnine_unit ninexnine_unit_122(
				.clk(clk),
				.rstn(rstn),
				.a0(P02C2),
				.a1(P02D2),
				.a2(P02E2),
				.a3(P03C2),
				.a4(P03D2),
				.a5(P03E2),
				.a6(P04C2),
				.a7(P04D2),
				.a8(P04E2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c022C0)
);

assign C02C0=c002C0+c012C0+c022C0;
assign A02C0=(C02C0>=0)?1:0;

ninexnine_unit ninexnine_unit_123(
				.clk(clk),
				.rstn(rstn),
				.a0(P02D0),
				.a1(P02E0),
				.a2(P02F0),
				.a3(P03D0),
				.a4(P03E0),
				.a5(P03F0),
				.a6(P04D0),
				.a7(P04E0),
				.a8(P04F0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c002D0)
);

ninexnine_unit ninexnine_unit_124(
				.clk(clk),
				.rstn(rstn),
				.a0(P02D1),
				.a1(P02E1),
				.a2(P02F1),
				.a3(P03D1),
				.a4(P03E1),
				.a5(P03F1),
				.a6(P04D1),
				.a7(P04E1),
				.a8(P04F1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c012D0)
);

ninexnine_unit ninexnine_unit_125(
				.clk(clk),
				.rstn(rstn),
				.a0(P02D2),
				.a1(P02E2),
				.a2(P02F2),
				.a3(P03D2),
				.a4(P03E2),
				.a5(P03F2),
				.a6(P04D2),
				.a7(P04E2),
				.a8(P04F2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c022D0)
);

assign C02D0=c002D0+c012D0+c022D0;
assign A02D0=(C02D0>=0)?1:0;

ninexnine_unit ninexnine_unit_126(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00300)
);

ninexnine_unit ninexnine_unit_127(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01300)
);

ninexnine_unit ninexnine_unit_128(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02300)
);

assign C0300=c00300+c01300+c02300;
assign A0300=(C0300>=0)?1:0;

ninexnine_unit ninexnine_unit_129(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00310)
);

ninexnine_unit ninexnine_unit_130(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01310)
);

ninexnine_unit ninexnine_unit_131(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02310)
);

assign C0310=c00310+c01310+c02310;
assign A0310=(C0310>=0)?1:0;

ninexnine_unit ninexnine_unit_132(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00320)
);

ninexnine_unit ninexnine_unit_133(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01320)
);

ninexnine_unit ninexnine_unit_134(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02320)
);

assign C0320=c00320+c01320+c02320;
assign A0320=(C0320>=0)?1:0;

ninexnine_unit ninexnine_unit_135(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00330)
);

ninexnine_unit ninexnine_unit_136(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01330)
);

ninexnine_unit ninexnine_unit_137(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02330)
);

assign C0330=c00330+c01330+c02330;
assign A0330=(C0330>=0)?1:0;

ninexnine_unit ninexnine_unit_138(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00340)
);

ninexnine_unit ninexnine_unit_139(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01340)
);

ninexnine_unit ninexnine_unit_140(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02340)
);

assign C0340=c00340+c01340+c02340;
assign A0340=(C0340>=0)?1:0;

ninexnine_unit ninexnine_unit_141(
				.clk(clk),
				.rstn(rstn),
				.a0(P0350),
				.a1(P0360),
				.a2(P0370),
				.a3(P0450),
				.a4(P0460),
				.a5(P0470),
				.a6(P0550),
				.a7(P0560),
				.a8(P0570),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00350)
);

ninexnine_unit ninexnine_unit_142(
				.clk(clk),
				.rstn(rstn),
				.a0(P0351),
				.a1(P0361),
				.a2(P0371),
				.a3(P0451),
				.a4(P0461),
				.a5(P0471),
				.a6(P0551),
				.a7(P0561),
				.a8(P0571),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01350)
);

ninexnine_unit ninexnine_unit_143(
				.clk(clk),
				.rstn(rstn),
				.a0(P0352),
				.a1(P0362),
				.a2(P0372),
				.a3(P0452),
				.a4(P0462),
				.a5(P0472),
				.a6(P0552),
				.a7(P0562),
				.a8(P0572),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02350)
);

assign C0350=c00350+c01350+c02350;
assign A0350=(C0350>=0)?1:0;

ninexnine_unit ninexnine_unit_144(
				.clk(clk),
				.rstn(rstn),
				.a0(P0360),
				.a1(P0370),
				.a2(P0380),
				.a3(P0460),
				.a4(P0470),
				.a5(P0480),
				.a6(P0560),
				.a7(P0570),
				.a8(P0580),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00360)
);

ninexnine_unit ninexnine_unit_145(
				.clk(clk),
				.rstn(rstn),
				.a0(P0361),
				.a1(P0371),
				.a2(P0381),
				.a3(P0461),
				.a4(P0471),
				.a5(P0481),
				.a6(P0561),
				.a7(P0571),
				.a8(P0581),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01360)
);

ninexnine_unit ninexnine_unit_146(
				.clk(clk),
				.rstn(rstn),
				.a0(P0362),
				.a1(P0372),
				.a2(P0382),
				.a3(P0462),
				.a4(P0472),
				.a5(P0482),
				.a6(P0562),
				.a7(P0572),
				.a8(P0582),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02360)
);

assign C0360=c00360+c01360+c02360;
assign A0360=(C0360>=0)?1:0;

ninexnine_unit ninexnine_unit_147(
				.clk(clk),
				.rstn(rstn),
				.a0(P0370),
				.a1(P0380),
				.a2(P0390),
				.a3(P0470),
				.a4(P0480),
				.a5(P0490),
				.a6(P0570),
				.a7(P0580),
				.a8(P0590),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00370)
);

ninexnine_unit ninexnine_unit_148(
				.clk(clk),
				.rstn(rstn),
				.a0(P0371),
				.a1(P0381),
				.a2(P0391),
				.a3(P0471),
				.a4(P0481),
				.a5(P0491),
				.a6(P0571),
				.a7(P0581),
				.a8(P0591),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01370)
);

ninexnine_unit ninexnine_unit_149(
				.clk(clk),
				.rstn(rstn),
				.a0(P0372),
				.a1(P0382),
				.a2(P0392),
				.a3(P0472),
				.a4(P0482),
				.a5(P0492),
				.a6(P0572),
				.a7(P0582),
				.a8(P0592),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02370)
);

assign C0370=c00370+c01370+c02370;
assign A0370=(C0370>=0)?1:0;

ninexnine_unit ninexnine_unit_150(
				.clk(clk),
				.rstn(rstn),
				.a0(P0380),
				.a1(P0390),
				.a2(P03A0),
				.a3(P0480),
				.a4(P0490),
				.a5(P04A0),
				.a6(P0580),
				.a7(P0590),
				.a8(P05A0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00380)
);

ninexnine_unit ninexnine_unit_151(
				.clk(clk),
				.rstn(rstn),
				.a0(P0381),
				.a1(P0391),
				.a2(P03A1),
				.a3(P0481),
				.a4(P0491),
				.a5(P04A1),
				.a6(P0581),
				.a7(P0591),
				.a8(P05A1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01380)
);

ninexnine_unit ninexnine_unit_152(
				.clk(clk),
				.rstn(rstn),
				.a0(P0382),
				.a1(P0392),
				.a2(P03A2),
				.a3(P0482),
				.a4(P0492),
				.a5(P04A2),
				.a6(P0582),
				.a7(P0592),
				.a8(P05A2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02380)
);

assign C0380=c00380+c01380+c02380;
assign A0380=(C0380>=0)?1:0;

ninexnine_unit ninexnine_unit_153(
				.clk(clk),
				.rstn(rstn),
				.a0(P0390),
				.a1(P03A0),
				.a2(P03B0),
				.a3(P0490),
				.a4(P04A0),
				.a5(P04B0),
				.a6(P0590),
				.a7(P05A0),
				.a8(P05B0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00390)
);

ninexnine_unit ninexnine_unit_154(
				.clk(clk),
				.rstn(rstn),
				.a0(P0391),
				.a1(P03A1),
				.a2(P03B1),
				.a3(P0491),
				.a4(P04A1),
				.a5(P04B1),
				.a6(P0591),
				.a7(P05A1),
				.a8(P05B1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01390)
);

ninexnine_unit ninexnine_unit_155(
				.clk(clk),
				.rstn(rstn),
				.a0(P0392),
				.a1(P03A2),
				.a2(P03B2),
				.a3(P0492),
				.a4(P04A2),
				.a5(P04B2),
				.a6(P0592),
				.a7(P05A2),
				.a8(P05B2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02390)
);

assign C0390=c00390+c01390+c02390;
assign A0390=(C0390>=0)?1:0;

ninexnine_unit ninexnine_unit_156(
				.clk(clk),
				.rstn(rstn),
				.a0(P03A0),
				.a1(P03B0),
				.a2(P03C0),
				.a3(P04A0),
				.a4(P04B0),
				.a5(P04C0),
				.a6(P05A0),
				.a7(P05B0),
				.a8(P05C0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c003A0)
);

ninexnine_unit ninexnine_unit_157(
				.clk(clk),
				.rstn(rstn),
				.a0(P03A1),
				.a1(P03B1),
				.a2(P03C1),
				.a3(P04A1),
				.a4(P04B1),
				.a5(P04C1),
				.a6(P05A1),
				.a7(P05B1),
				.a8(P05C1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c013A0)
);

ninexnine_unit ninexnine_unit_158(
				.clk(clk),
				.rstn(rstn),
				.a0(P03A2),
				.a1(P03B2),
				.a2(P03C2),
				.a3(P04A2),
				.a4(P04B2),
				.a5(P04C2),
				.a6(P05A2),
				.a7(P05B2),
				.a8(P05C2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c023A0)
);

assign C03A0=c003A0+c013A0+c023A0;
assign A03A0=(C03A0>=0)?1:0;

ninexnine_unit ninexnine_unit_159(
				.clk(clk),
				.rstn(rstn),
				.a0(P03B0),
				.a1(P03C0),
				.a2(P03D0),
				.a3(P04B0),
				.a4(P04C0),
				.a5(P04D0),
				.a6(P05B0),
				.a7(P05C0),
				.a8(P05D0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c003B0)
);

ninexnine_unit ninexnine_unit_160(
				.clk(clk),
				.rstn(rstn),
				.a0(P03B1),
				.a1(P03C1),
				.a2(P03D1),
				.a3(P04B1),
				.a4(P04C1),
				.a5(P04D1),
				.a6(P05B1),
				.a7(P05C1),
				.a8(P05D1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c013B0)
);

ninexnine_unit ninexnine_unit_161(
				.clk(clk),
				.rstn(rstn),
				.a0(P03B2),
				.a1(P03C2),
				.a2(P03D2),
				.a3(P04B2),
				.a4(P04C2),
				.a5(P04D2),
				.a6(P05B2),
				.a7(P05C2),
				.a8(P05D2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c023B0)
);

assign C03B0=c003B0+c013B0+c023B0;
assign A03B0=(C03B0>=0)?1:0;

ninexnine_unit ninexnine_unit_162(
				.clk(clk),
				.rstn(rstn),
				.a0(P03C0),
				.a1(P03D0),
				.a2(P03E0),
				.a3(P04C0),
				.a4(P04D0),
				.a5(P04E0),
				.a6(P05C0),
				.a7(P05D0),
				.a8(P05E0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c003C0)
);

ninexnine_unit ninexnine_unit_163(
				.clk(clk),
				.rstn(rstn),
				.a0(P03C1),
				.a1(P03D1),
				.a2(P03E1),
				.a3(P04C1),
				.a4(P04D1),
				.a5(P04E1),
				.a6(P05C1),
				.a7(P05D1),
				.a8(P05E1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c013C0)
);

ninexnine_unit ninexnine_unit_164(
				.clk(clk),
				.rstn(rstn),
				.a0(P03C2),
				.a1(P03D2),
				.a2(P03E2),
				.a3(P04C2),
				.a4(P04D2),
				.a5(P04E2),
				.a6(P05C2),
				.a7(P05D2),
				.a8(P05E2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c023C0)
);

assign C03C0=c003C0+c013C0+c023C0;
assign A03C0=(C03C0>=0)?1:0;

ninexnine_unit ninexnine_unit_165(
				.clk(clk),
				.rstn(rstn),
				.a0(P03D0),
				.a1(P03E0),
				.a2(P03F0),
				.a3(P04D0),
				.a4(P04E0),
				.a5(P04F0),
				.a6(P05D0),
				.a7(P05E0),
				.a8(P05F0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c003D0)
);

ninexnine_unit ninexnine_unit_166(
				.clk(clk),
				.rstn(rstn),
				.a0(P03D1),
				.a1(P03E1),
				.a2(P03F1),
				.a3(P04D1),
				.a4(P04E1),
				.a5(P04F1),
				.a6(P05D1),
				.a7(P05E1),
				.a8(P05F1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c013D0)
);

ninexnine_unit ninexnine_unit_167(
				.clk(clk),
				.rstn(rstn),
				.a0(P03D2),
				.a1(P03E2),
				.a2(P03F2),
				.a3(P04D2),
				.a4(P04E2),
				.a5(P04F2),
				.a6(P05D2),
				.a7(P05E2),
				.a8(P05F2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c023D0)
);

assign C03D0=c003D0+c013D0+c023D0;
assign A03D0=(C03D0>=0)?1:0;

ninexnine_unit ninexnine_unit_168(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00400)
);

ninexnine_unit ninexnine_unit_169(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01400)
);

ninexnine_unit ninexnine_unit_170(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02400)
);

assign C0400=c00400+c01400+c02400;
assign A0400=(C0400>=0)?1:0;

ninexnine_unit ninexnine_unit_171(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00410)
);

ninexnine_unit ninexnine_unit_172(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01410)
);

ninexnine_unit ninexnine_unit_173(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02410)
);

assign C0410=c00410+c01410+c02410;
assign A0410=(C0410>=0)?1:0;

ninexnine_unit ninexnine_unit_174(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00420)
);

ninexnine_unit ninexnine_unit_175(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01420)
);

ninexnine_unit ninexnine_unit_176(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02420)
);

assign C0420=c00420+c01420+c02420;
assign A0420=(C0420>=0)?1:0;

ninexnine_unit ninexnine_unit_177(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00430)
);

ninexnine_unit ninexnine_unit_178(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01430)
);

ninexnine_unit ninexnine_unit_179(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02430)
);

assign C0430=c00430+c01430+c02430;
assign A0430=(C0430>=0)?1:0;

ninexnine_unit ninexnine_unit_180(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00440)
);

ninexnine_unit ninexnine_unit_181(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01440)
);

ninexnine_unit ninexnine_unit_182(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02440)
);

assign C0440=c00440+c01440+c02440;
assign A0440=(C0440>=0)?1:0;

ninexnine_unit ninexnine_unit_183(
				.clk(clk),
				.rstn(rstn),
				.a0(P0450),
				.a1(P0460),
				.a2(P0470),
				.a3(P0550),
				.a4(P0560),
				.a5(P0570),
				.a6(P0650),
				.a7(P0660),
				.a8(P0670),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00450)
);

ninexnine_unit ninexnine_unit_184(
				.clk(clk),
				.rstn(rstn),
				.a0(P0451),
				.a1(P0461),
				.a2(P0471),
				.a3(P0551),
				.a4(P0561),
				.a5(P0571),
				.a6(P0651),
				.a7(P0661),
				.a8(P0671),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01450)
);

ninexnine_unit ninexnine_unit_185(
				.clk(clk),
				.rstn(rstn),
				.a0(P0452),
				.a1(P0462),
				.a2(P0472),
				.a3(P0552),
				.a4(P0562),
				.a5(P0572),
				.a6(P0652),
				.a7(P0662),
				.a8(P0672),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02450)
);

assign C0450=c00450+c01450+c02450;
assign A0450=(C0450>=0)?1:0;

ninexnine_unit ninexnine_unit_186(
				.clk(clk),
				.rstn(rstn),
				.a0(P0460),
				.a1(P0470),
				.a2(P0480),
				.a3(P0560),
				.a4(P0570),
				.a5(P0580),
				.a6(P0660),
				.a7(P0670),
				.a8(P0680),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00460)
);

ninexnine_unit ninexnine_unit_187(
				.clk(clk),
				.rstn(rstn),
				.a0(P0461),
				.a1(P0471),
				.a2(P0481),
				.a3(P0561),
				.a4(P0571),
				.a5(P0581),
				.a6(P0661),
				.a7(P0671),
				.a8(P0681),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01460)
);

ninexnine_unit ninexnine_unit_188(
				.clk(clk),
				.rstn(rstn),
				.a0(P0462),
				.a1(P0472),
				.a2(P0482),
				.a3(P0562),
				.a4(P0572),
				.a5(P0582),
				.a6(P0662),
				.a7(P0672),
				.a8(P0682),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02460)
);

assign C0460=c00460+c01460+c02460;
assign A0460=(C0460>=0)?1:0;

ninexnine_unit ninexnine_unit_189(
				.clk(clk),
				.rstn(rstn),
				.a0(P0470),
				.a1(P0480),
				.a2(P0490),
				.a3(P0570),
				.a4(P0580),
				.a5(P0590),
				.a6(P0670),
				.a7(P0680),
				.a8(P0690),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00470)
);

ninexnine_unit ninexnine_unit_190(
				.clk(clk),
				.rstn(rstn),
				.a0(P0471),
				.a1(P0481),
				.a2(P0491),
				.a3(P0571),
				.a4(P0581),
				.a5(P0591),
				.a6(P0671),
				.a7(P0681),
				.a8(P0691),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01470)
);

ninexnine_unit ninexnine_unit_191(
				.clk(clk),
				.rstn(rstn),
				.a0(P0472),
				.a1(P0482),
				.a2(P0492),
				.a3(P0572),
				.a4(P0582),
				.a5(P0592),
				.a6(P0672),
				.a7(P0682),
				.a8(P0692),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02470)
);

assign C0470=c00470+c01470+c02470;
assign A0470=(C0470>=0)?1:0;

ninexnine_unit ninexnine_unit_192(
				.clk(clk),
				.rstn(rstn),
				.a0(P0480),
				.a1(P0490),
				.a2(P04A0),
				.a3(P0580),
				.a4(P0590),
				.a5(P05A0),
				.a6(P0680),
				.a7(P0690),
				.a8(P06A0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00480)
);

ninexnine_unit ninexnine_unit_193(
				.clk(clk),
				.rstn(rstn),
				.a0(P0481),
				.a1(P0491),
				.a2(P04A1),
				.a3(P0581),
				.a4(P0591),
				.a5(P05A1),
				.a6(P0681),
				.a7(P0691),
				.a8(P06A1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01480)
);

ninexnine_unit ninexnine_unit_194(
				.clk(clk),
				.rstn(rstn),
				.a0(P0482),
				.a1(P0492),
				.a2(P04A2),
				.a3(P0582),
				.a4(P0592),
				.a5(P05A2),
				.a6(P0682),
				.a7(P0692),
				.a8(P06A2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02480)
);

assign C0480=c00480+c01480+c02480;
assign A0480=(C0480>=0)?1:0;

ninexnine_unit ninexnine_unit_195(
				.clk(clk),
				.rstn(rstn),
				.a0(P0490),
				.a1(P04A0),
				.a2(P04B0),
				.a3(P0590),
				.a4(P05A0),
				.a5(P05B0),
				.a6(P0690),
				.a7(P06A0),
				.a8(P06B0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00490)
);

ninexnine_unit ninexnine_unit_196(
				.clk(clk),
				.rstn(rstn),
				.a0(P0491),
				.a1(P04A1),
				.a2(P04B1),
				.a3(P0591),
				.a4(P05A1),
				.a5(P05B1),
				.a6(P0691),
				.a7(P06A1),
				.a8(P06B1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01490)
);

ninexnine_unit ninexnine_unit_197(
				.clk(clk),
				.rstn(rstn),
				.a0(P0492),
				.a1(P04A2),
				.a2(P04B2),
				.a3(P0592),
				.a4(P05A2),
				.a5(P05B2),
				.a6(P0692),
				.a7(P06A2),
				.a8(P06B2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02490)
);

assign C0490=c00490+c01490+c02490;
assign A0490=(C0490>=0)?1:0;

ninexnine_unit ninexnine_unit_198(
				.clk(clk),
				.rstn(rstn),
				.a0(P04A0),
				.a1(P04B0),
				.a2(P04C0),
				.a3(P05A0),
				.a4(P05B0),
				.a5(P05C0),
				.a6(P06A0),
				.a7(P06B0),
				.a8(P06C0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c004A0)
);

ninexnine_unit ninexnine_unit_199(
				.clk(clk),
				.rstn(rstn),
				.a0(P04A1),
				.a1(P04B1),
				.a2(P04C1),
				.a3(P05A1),
				.a4(P05B1),
				.a5(P05C1),
				.a6(P06A1),
				.a7(P06B1),
				.a8(P06C1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c014A0)
);

ninexnine_unit ninexnine_unit_200(
				.clk(clk),
				.rstn(rstn),
				.a0(P04A2),
				.a1(P04B2),
				.a2(P04C2),
				.a3(P05A2),
				.a4(P05B2),
				.a5(P05C2),
				.a6(P06A2),
				.a7(P06B2),
				.a8(P06C2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c024A0)
);

assign C04A0=c004A0+c014A0+c024A0;
assign A04A0=(C04A0>=0)?1:0;

ninexnine_unit ninexnine_unit_201(
				.clk(clk),
				.rstn(rstn),
				.a0(P04B0),
				.a1(P04C0),
				.a2(P04D0),
				.a3(P05B0),
				.a4(P05C0),
				.a5(P05D0),
				.a6(P06B0),
				.a7(P06C0),
				.a8(P06D0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c004B0)
);

ninexnine_unit ninexnine_unit_202(
				.clk(clk),
				.rstn(rstn),
				.a0(P04B1),
				.a1(P04C1),
				.a2(P04D1),
				.a3(P05B1),
				.a4(P05C1),
				.a5(P05D1),
				.a6(P06B1),
				.a7(P06C1),
				.a8(P06D1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c014B0)
);

ninexnine_unit ninexnine_unit_203(
				.clk(clk),
				.rstn(rstn),
				.a0(P04B2),
				.a1(P04C2),
				.a2(P04D2),
				.a3(P05B2),
				.a4(P05C2),
				.a5(P05D2),
				.a6(P06B2),
				.a7(P06C2),
				.a8(P06D2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c024B0)
);

assign C04B0=c004B0+c014B0+c024B0;
assign A04B0=(C04B0>=0)?1:0;

ninexnine_unit ninexnine_unit_204(
				.clk(clk),
				.rstn(rstn),
				.a0(P04C0),
				.a1(P04D0),
				.a2(P04E0),
				.a3(P05C0),
				.a4(P05D0),
				.a5(P05E0),
				.a6(P06C0),
				.a7(P06D0),
				.a8(P06E0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c004C0)
);

ninexnine_unit ninexnine_unit_205(
				.clk(clk),
				.rstn(rstn),
				.a0(P04C1),
				.a1(P04D1),
				.a2(P04E1),
				.a3(P05C1),
				.a4(P05D1),
				.a5(P05E1),
				.a6(P06C1),
				.a7(P06D1),
				.a8(P06E1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c014C0)
);

ninexnine_unit ninexnine_unit_206(
				.clk(clk),
				.rstn(rstn),
				.a0(P04C2),
				.a1(P04D2),
				.a2(P04E2),
				.a3(P05C2),
				.a4(P05D2),
				.a5(P05E2),
				.a6(P06C2),
				.a7(P06D2),
				.a8(P06E2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c024C0)
);

assign C04C0=c004C0+c014C0+c024C0;
assign A04C0=(C04C0>=0)?1:0;

ninexnine_unit ninexnine_unit_207(
				.clk(clk),
				.rstn(rstn),
				.a0(P04D0),
				.a1(P04E0),
				.a2(P04F0),
				.a3(P05D0),
				.a4(P05E0),
				.a5(P05F0),
				.a6(P06D0),
				.a7(P06E0),
				.a8(P06F0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c004D0)
);

ninexnine_unit ninexnine_unit_208(
				.clk(clk),
				.rstn(rstn),
				.a0(P04D1),
				.a1(P04E1),
				.a2(P04F1),
				.a3(P05D1),
				.a4(P05E1),
				.a5(P05F1),
				.a6(P06D1),
				.a7(P06E1),
				.a8(P06F1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c014D0)
);

ninexnine_unit ninexnine_unit_209(
				.clk(clk),
				.rstn(rstn),
				.a0(P04D2),
				.a1(P04E2),
				.a2(P04F2),
				.a3(P05D2),
				.a4(P05E2),
				.a5(P05F2),
				.a6(P06D2),
				.a7(P06E2),
				.a8(P06F2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c024D0)
);

assign C04D0=c004D0+c014D0+c024D0;
assign A04D0=(C04D0>=0)?1:0;

ninexnine_unit ninexnine_unit_210(
				.clk(clk),
				.rstn(rstn),
				.a0(P0500),
				.a1(P0510),
				.a2(P0520),
				.a3(P0600),
				.a4(P0610),
				.a5(P0620),
				.a6(P0700),
				.a7(P0710),
				.a8(P0720),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00500)
);

ninexnine_unit ninexnine_unit_211(
				.clk(clk),
				.rstn(rstn),
				.a0(P0501),
				.a1(P0511),
				.a2(P0521),
				.a3(P0601),
				.a4(P0611),
				.a5(P0621),
				.a6(P0701),
				.a7(P0711),
				.a8(P0721),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01500)
);

ninexnine_unit ninexnine_unit_212(
				.clk(clk),
				.rstn(rstn),
				.a0(P0502),
				.a1(P0512),
				.a2(P0522),
				.a3(P0602),
				.a4(P0612),
				.a5(P0622),
				.a6(P0702),
				.a7(P0712),
				.a8(P0722),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02500)
);

assign C0500=c00500+c01500+c02500;
assign A0500=(C0500>=0)?1:0;

ninexnine_unit ninexnine_unit_213(
				.clk(clk),
				.rstn(rstn),
				.a0(P0510),
				.a1(P0520),
				.a2(P0530),
				.a3(P0610),
				.a4(P0620),
				.a5(P0630),
				.a6(P0710),
				.a7(P0720),
				.a8(P0730),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00510)
);

ninexnine_unit ninexnine_unit_214(
				.clk(clk),
				.rstn(rstn),
				.a0(P0511),
				.a1(P0521),
				.a2(P0531),
				.a3(P0611),
				.a4(P0621),
				.a5(P0631),
				.a6(P0711),
				.a7(P0721),
				.a8(P0731),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01510)
);

ninexnine_unit ninexnine_unit_215(
				.clk(clk),
				.rstn(rstn),
				.a0(P0512),
				.a1(P0522),
				.a2(P0532),
				.a3(P0612),
				.a4(P0622),
				.a5(P0632),
				.a6(P0712),
				.a7(P0722),
				.a8(P0732),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02510)
);

assign C0510=c00510+c01510+c02510;
assign A0510=(C0510>=0)?1:0;

ninexnine_unit ninexnine_unit_216(
				.clk(clk),
				.rstn(rstn),
				.a0(P0520),
				.a1(P0530),
				.a2(P0540),
				.a3(P0620),
				.a4(P0630),
				.a5(P0640),
				.a6(P0720),
				.a7(P0730),
				.a8(P0740),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00520)
);

ninexnine_unit ninexnine_unit_217(
				.clk(clk),
				.rstn(rstn),
				.a0(P0521),
				.a1(P0531),
				.a2(P0541),
				.a3(P0621),
				.a4(P0631),
				.a5(P0641),
				.a6(P0721),
				.a7(P0731),
				.a8(P0741),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01520)
);

ninexnine_unit ninexnine_unit_218(
				.clk(clk),
				.rstn(rstn),
				.a0(P0522),
				.a1(P0532),
				.a2(P0542),
				.a3(P0622),
				.a4(P0632),
				.a5(P0642),
				.a6(P0722),
				.a7(P0732),
				.a8(P0742),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02520)
);

assign C0520=c00520+c01520+c02520;
assign A0520=(C0520>=0)?1:0;

ninexnine_unit ninexnine_unit_219(
				.clk(clk),
				.rstn(rstn),
				.a0(P0530),
				.a1(P0540),
				.a2(P0550),
				.a3(P0630),
				.a4(P0640),
				.a5(P0650),
				.a6(P0730),
				.a7(P0740),
				.a8(P0750),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00530)
);

ninexnine_unit ninexnine_unit_220(
				.clk(clk),
				.rstn(rstn),
				.a0(P0531),
				.a1(P0541),
				.a2(P0551),
				.a3(P0631),
				.a4(P0641),
				.a5(P0651),
				.a6(P0731),
				.a7(P0741),
				.a8(P0751),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01530)
);

ninexnine_unit ninexnine_unit_221(
				.clk(clk),
				.rstn(rstn),
				.a0(P0532),
				.a1(P0542),
				.a2(P0552),
				.a3(P0632),
				.a4(P0642),
				.a5(P0652),
				.a6(P0732),
				.a7(P0742),
				.a8(P0752),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02530)
);

assign C0530=c00530+c01530+c02530;
assign A0530=(C0530>=0)?1:0;

ninexnine_unit ninexnine_unit_222(
				.clk(clk),
				.rstn(rstn),
				.a0(P0540),
				.a1(P0550),
				.a2(P0560),
				.a3(P0640),
				.a4(P0650),
				.a5(P0660),
				.a6(P0740),
				.a7(P0750),
				.a8(P0760),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00540)
);

ninexnine_unit ninexnine_unit_223(
				.clk(clk),
				.rstn(rstn),
				.a0(P0541),
				.a1(P0551),
				.a2(P0561),
				.a3(P0641),
				.a4(P0651),
				.a5(P0661),
				.a6(P0741),
				.a7(P0751),
				.a8(P0761),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01540)
);

ninexnine_unit ninexnine_unit_224(
				.clk(clk),
				.rstn(rstn),
				.a0(P0542),
				.a1(P0552),
				.a2(P0562),
				.a3(P0642),
				.a4(P0652),
				.a5(P0662),
				.a6(P0742),
				.a7(P0752),
				.a8(P0762),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02540)
);

assign C0540=c00540+c01540+c02540;
assign A0540=(C0540>=0)?1:0;

ninexnine_unit ninexnine_unit_225(
				.clk(clk),
				.rstn(rstn),
				.a0(P0550),
				.a1(P0560),
				.a2(P0570),
				.a3(P0650),
				.a4(P0660),
				.a5(P0670),
				.a6(P0750),
				.a7(P0760),
				.a8(P0770),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00550)
);

ninexnine_unit ninexnine_unit_226(
				.clk(clk),
				.rstn(rstn),
				.a0(P0551),
				.a1(P0561),
				.a2(P0571),
				.a3(P0651),
				.a4(P0661),
				.a5(P0671),
				.a6(P0751),
				.a7(P0761),
				.a8(P0771),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01550)
);

ninexnine_unit ninexnine_unit_227(
				.clk(clk),
				.rstn(rstn),
				.a0(P0552),
				.a1(P0562),
				.a2(P0572),
				.a3(P0652),
				.a4(P0662),
				.a5(P0672),
				.a6(P0752),
				.a7(P0762),
				.a8(P0772),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02550)
);

assign C0550=c00550+c01550+c02550;
assign A0550=(C0550>=0)?1:0;

ninexnine_unit ninexnine_unit_228(
				.clk(clk),
				.rstn(rstn),
				.a0(P0560),
				.a1(P0570),
				.a2(P0580),
				.a3(P0660),
				.a4(P0670),
				.a5(P0680),
				.a6(P0760),
				.a7(P0770),
				.a8(P0780),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00560)
);

ninexnine_unit ninexnine_unit_229(
				.clk(clk),
				.rstn(rstn),
				.a0(P0561),
				.a1(P0571),
				.a2(P0581),
				.a3(P0661),
				.a4(P0671),
				.a5(P0681),
				.a6(P0761),
				.a7(P0771),
				.a8(P0781),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01560)
);

ninexnine_unit ninexnine_unit_230(
				.clk(clk),
				.rstn(rstn),
				.a0(P0562),
				.a1(P0572),
				.a2(P0582),
				.a3(P0662),
				.a4(P0672),
				.a5(P0682),
				.a6(P0762),
				.a7(P0772),
				.a8(P0782),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02560)
);

assign C0560=c00560+c01560+c02560;
assign A0560=(C0560>=0)?1:0;

ninexnine_unit ninexnine_unit_231(
				.clk(clk),
				.rstn(rstn),
				.a0(P0570),
				.a1(P0580),
				.a2(P0590),
				.a3(P0670),
				.a4(P0680),
				.a5(P0690),
				.a6(P0770),
				.a7(P0780),
				.a8(P0790),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00570)
);

ninexnine_unit ninexnine_unit_232(
				.clk(clk),
				.rstn(rstn),
				.a0(P0571),
				.a1(P0581),
				.a2(P0591),
				.a3(P0671),
				.a4(P0681),
				.a5(P0691),
				.a6(P0771),
				.a7(P0781),
				.a8(P0791),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01570)
);

ninexnine_unit ninexnine_unit_233(
				.clk(clk),
				.rstn(rstn),
				.a0(P0572),
				.a1(P0582),
				.a2(P0592),
				.a3(P0672),
				.a4(P0682),
				.a5(P0692),
				.a6(P0772),
				.a7(P0782),
				.a8(P0792),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02570)
);

assign C0570=c00570+c01570+c02570;
assign A0570=(C0570>=0)?1:0;

ninexnine_unit ninexnine_unit_234(
				.clk(clk),
				.rstn(rstn),
				.a0(P0580),
				.a1(P0590),
				.a2(P05A0),
				.a3(P0680),
				.a4(P0690),
				.a5(P06A0),
				.a6(P0780),
				.a7(P0790),
				.a8(P07A0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00580)
);

ninexnine_unit ninexnine_unit_235(
				.clk(clk),
				.rstn(rstn),
				.a0(P0581),
				.a1(P0591),
				.a2(P05A1),
				.a3(P0681),
				.a4(P0691),
				.a5(P06A1),
				.a6(P0781),
				.a7(P0791),
				.a8(P07A1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01580)
);

ninexnine_unit ninexnine_unit_236(
				.clk(clk),
				.rstn(rstn),
				.a0(P0582),
				.a1(P0592),
				.a2(P05A2),
				.a3(P0682),
				.a4(P0692),
				.a5(P06A2),
				.a6(P0782),
				.a7(P0792),
				.a8(P07A2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02580)
);

assign C0580=c00580+c01580+c02580;
assign A0580=(C0580>=0)?1:0;

ninexnine_unit ninexnine_unit_237(
				.clk(clk),
				.rstn(rstn),
				.a0(P0590),
				.a1(P05A0),
				.a2(P05B0),
				.a3(P0690),
				.a4(P06A0),
				.a5(P06B0),
				.a6(P0790),
				.a7(P07A0),
				.a8(P07B0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00590)
);

ninexnine_unit ninexnine_unit_238(
				.clk(clk),
				.rstn(rstn),
				.a0(P0591),
				.a1(P05A1),
				.a2(P05B1),
				.a3(P0691),
				.a4(P06A1),
				.a5(P06B1),
				.a6(P0791),
				.a7(P07A1),
				.a8(P07B1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01590)
);

ninexnine_unit ninexnine_unit_239(
				.clk(clk),
				.rstn(rstn),
				.a0(P0592),
				.a1(P05A2),
				.a2(P05B2),
				.a3(P0692),
				.a4(P06A2),
				.a5(P06B2),
				.a6(P0792),
				.a7(P07A2),
				.a8(P07B2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02590)
);

assign C0590=c00590+c01590+c02590;
assign A0590=(C0590>=0)?1:0;

ninexnine_unit ninexnine_unit_240(
				.clk(clk),
				.rstn(rstn),
				.a0(P05A0),
				.a1(P05B0),
				.a2(P05C0),
				.a3(P06A0),
				.a4(P06B0),
				.a5(P06C0),
				.a6(P07A0),
				.a7(P07B0),
				.a8(P07C0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c005A0)
);

ninexnine_unit ninexnine_unit_241(
				.clk(clk),
				.rstn(rstn),
				.a0(P05A1),
				.a1(P05B1),
				.a2(P05C1),
				.a3(P06A1),
				.a4(P06B1),
				.a5(P06C1),
				.a6(P07A1),
				.a7(P07B1),
				.a8(P07C1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c015A0)
);

ninexnine_unit ninexnine_unit_242(
				.clk(clk),
				.rstn(rstn),
				.a0(P05A2),
				.a1(P05B2),
				.a2(P05C2),
				.a3(P06A2),
				.a4(P06B2),
				.a5(P06C2),
				.a6(P07A2),
				.a7(P07B2),
				.a8(P07C2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c025A0)
);

assign C05A0=c005A0+c015A0+c025A0;
assign A05A0=(C05A0>=0)?1:0;

ninexnine_unit ninexnine_unit_243(
				.clk(clk),
				.rstn(rstn),
				.a0(P05B0),
				.a1(P05C0),
				.a2(P05D0),
				.a3(P06B0),
				.a4(P06C0),
				.a5(P06D0),
				.a6(P07B0),
				.a7(P07C0),
				.a8(P07D0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c005B0)
);

ninexnine_unit ninexnine_unit_244(
				.clk(clk),
				.rstn(rstn),
				.a0(P05B1),
				.a1(P05C1),
				.a2(P05D1),
				.a3(P06B1),
				.a4(P06C1),
				.a5(P06D1),
				.a6(P07B1),
				.a7(P07C1),
				.a8(P07D1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c015B0)
);

ninexnine_unit ninexnine_unit_245(
				.clk(clk),
				.rstn(rstn),
				.a0(P05B2),
				.a1(P05C2),
				.a2(P05D2),
				.a3(P06B2),
				.a4(P06C2),
				.a5(P06D2),
				.a6(P07B2),
				.a7(P07C2),
				.a8(P07D2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c025B0)
);

assign C05B0=c005B0+c015B0+c025B0;
assign A05B0=(C05B0>=0)?1:0;

ninexnine_unit ninexnine_unit_246(
				.clk(clk),
				.rstn(rstn),
				.a0(P05C0),
				.a1(P05D0),
				.a2(P05E0),
				.a3(P06C0),
				.a4(P06D0),
				.a5(P06E0),
				.a6(P07C0),
				.a7(P07D0),
				.a8(P07E0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c005C0)
);

ninexnine_unit ninexnine_unit_247(
				.clk(clk),
				.rstn(rstn),
				.a0(P05C1),
				.a1(P05D1),
				.a2(P05E1),
				.a3(P06C1),
				.a4(P06D1),
				.a5(P06E1),
				.a6(P07C1),
				.a7(P07D1),
				.a8(P07E1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c015C0)
);

ninexnine_unit ninexnine_unit_248(
				.clk(clk),
				.rstn(rstn),
				.a0(P05C2),
				.a1(P05D2),
				.a2(P05E2),
				.a3(P06C2),
				.a4(P06D2),
				.a5(P06E2),
				.a6(P07C2),
				.a7(P07D2),
				.a8(P07E2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c025C0)
);

assign C05C0=c005C0+c015C0+c025C0;
assign A05C0=(C05C0>=0)?1:0;

ninexnine_unit ninexnine_unit_249(
				.clk(clk),
				.rstn(rstn),
				.a0(P05D0),
				.a1(P05E0),
				.a2(P05F0),
				.a3(P06D0),
				.a4(P06E0),
				.a5(P06F0),
				.a6(P07D0),
				.a7(P07E0),
				.a8(P07F0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c005D0)
);

ninexnine_unit ninexnine_unit_250(
				.clk(clk),
				.rstn(rstn),
				.a0(P05D1),
				.a1(P05E1),
				.a2(P05F1),
				.a3(P06D1),
				.a4(P06E1),
				.a5(P06F1),
				.a6(P07D1),
				.a7(P07E1),
				.a8(P07F1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c015D0)
);

ninexnine_unit ninexnine_unit_251(
				.clk(clk),
				.rstn(rstn),
				.a0(P05D2),
				.a1(P05E2),
				.a2(P05F2),
				.a3(P06D2),
				.a4(P06E2),
				.a5(P06F2),
				.a6(P07D2),
				.a7(P07E2),
				.a8(P07F2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c025D0)
);

assign C05D0=c005D0+c015D0+c025D0;
assign A05D0=(C05D0>=0)?1:0;

ninexnine_unit ninexnine_unit_252(
				.clk(clk),
				.rstn(rstn),
				.a0(P0600),
				.a1(P0610),
				.a2(P0620),
				.a3(P0700),
				.a4(P0710),
				.a5(P0720),
				.a6(P0800),
				.a7(P0810),
				.a8(P0820),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00600)
);

ninexnine_unit ninexnine_unit_253(
				.clk(clk),
				.rstn(rstn),
				.a0(P0601),
				.a1(P0611),
				.a2(P0621),
				.a3(P0701),
				.a4(P0711),
				.a5(P0721),
				.a6(P0801),
				.a7(P0811),
				.a8(P0821),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01600)
);

ninexnine_unit ninexnine_unit_254(
				.clk(clk),
				.rstn(rstn),
				.a0(P0602),
				.a1(P0612),
				.a2(P0622),
				.a3(P0702),
				.a4(P0712),
				.a5(P0722),
				.a6(P0802),
				.a7(P0812),
				.a8(P0822),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02600)
);

assign C0600=c00600+c01600+c02600;
assign A0600=(C0600>=0)?1:0;

ninexnine_unit ninexnine_unit_255(
				.clk(clk),
				.rstn(rstn),
				.a0(P0610),
				.a1(P0620),
				.a2(P0630),
				.a3(P0710),
				.a4(P0720),
				.a5(P0730),
				.a6(P0810),
				.a7(P0820),
				.a8(P0830),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00610)
);

ninexnine_unit ninexnine_unit_256(
				.clk(clk),
				.rstn(rstn),
				.a0(P0611),
				.a1(P0621),
				.a2(P0631),
				.a3(P0711),
				.a4(P0721),
				.a5(P0731),
				.a6(P0811),
				.a7(P0821),
				.a8(P0831),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01610)
);

ninexnine_unit ninexnine_unit_257(
				.clk(clk),
				.rstn(rstn),
				.a0(P0612),
				.a1(P0622),
				.a2(P0632),
				.a3(P0712),
				.a4(P0722),
				.a5(P0732),
				.a6(P0812),
				.a7(P0822),
				.a8(P0832),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02610)
);

assign C0610=c00610+c01610+c02610;
assign A0610=(C0610>=0)?1:0;

ninexnine_unit ninexnine_unit_258(
				.clk(clk),
				.rstn(rstn),
				.a0(P0620),
				.a1(P0630),
				.a2(P0640),
				.a3(P0720),
				.a4(P0730),
				.a5(P0740),
				.a6(P0820),
				.a7(P0830),
				.a8(P0840),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00620)
);

ninexnine_unit ninexnine_unit_259(
				.clk(clk),
				.rstn(rstn),
				.a0(P0621),
				.a1(P0631),
				.a2(P0641),
				.a3(P0721),
				.a4(P0731),
				.a5(P0741),
				.a6(P0821),
				.a7(P0831),
				.a8(P0841),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01620)
);

ninexnine_unit ninexnine_unit_260(
				.clk(clk),
				.rstn(rstn),
				.a0(P0622),
				.a1(P0632),
				.a2(P0642),
				.a3(P0722),
				.a4(P0732),
				.a5(P0742),
				.a6(P0822),
				.a7(P0832),
				.a8(P0842),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02620)
);

assign C0620=c00620+c01620+c02620;
assign A0620=(C0620>=0)?1:0;

ninexnine_unit ninexnine_unit_261(
				.clk(clk),
				.rstn(rstn),
				.a0(P0630),
				.a1(P0640),
				.a2(P0650),
				.a3(P0730),
				.a4(P0740),
				.a5(P0750),
				.a6(P0830),
				.a7(P0840),
				.a8(P0850),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00630)
);

ninexnine_unit ninexnine_unit_262(
				.clk(clk),
				.rstn(rstn),
				.a0(P0631),
				.a1(P0641),
				.a2(P0651),
				.a3(P0731),
				.a4(P0741),
				.a5(P0751),
				.a6(P0831),
				.a7(P0841),
				.a8(P0851),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01630)
);

ninexnine_unit ninexnine_unit_263(
				.clk(clk),
				.rstn(rstn),
				.a0(P0632),
				.a1(P0642),
				.a2(P0652),
				.a3(P0732),
				.a4(P0742),
				.a5(P0752),
				.a6(P0832),
				.a7(P0842),
				.a8(P0852),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02630)
);

assign C0630=c00630+c01630+c02630;
assign A0630=(C0630>=0)?1:0;

ninexnine_unit ninexnine_unit_264(
				.clk(clk),
				.rstn(rstn),
				.a0(P0640),
				.a1(P0650),
				.a2(P0660),
				.a3(P0740),
				.a4(P0750),
				.a5(P0760),
				.a6(P0840),
				.a7(P0850),
				.a8(P0860),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00640)
);

ninexnine_unit ninexnine_unit_265(
				.clk(clk),
				.rstn(rstn),
				.a0(P0641),
				.a1(P0651),
				.a2(P0661),
				.a3(P0741),
				.a4(P0751),
				.a5(P0761),
				.a6(P0841),
				.a7(P0851),
				.a8(P0861),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01640)
);

ninexnine_unit ninexnine_unit_266(
				.clk(clk),
				.rstn(rstn),
				.a0(P0642),
				.a1(P0652),
				.a2(P0662),
				.a3(P0742),
				.a4(P0752),
				.a5(P0762),
				.a6(P0842),
				.a7(P0852),
				.a8(P0862),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02640)
);

assign C0640=c00640+c01640+c02640;
assign A0640=(C0640>=0)?1:0;

ninexnine_unit ninexnine_unit_267(
				.clk(clk),
				.rstn(rstn),
				.a0(P0650),
				.a1(P0660),
				.a2(P0670),
				.a3(P0750),
				.a4(P0760),
				.a5(P0770),
				.a6(P0850),
				.a7(P0860),
				.a8(P0870),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00650)
);

ninexnine_unit ninexnine_unit_268(
				.clk(clk),
				.rstn(rstn),
				.a0(P0651),
				.a1(P0661),
				.a2(P0671),
				.a3(P0751),
				.a4(P0761),
				.a5(P0771),
				.a6(P0851),
				.a7(P0861),
				.a8(P0871),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01650)
);

ninexnine_unit ninexnine_unit_269(
				.clk(clk),
				.rstn(rstn),
				.a0(P0652),
				.a1(P0662),
				.a2(P0672),
				.a3(P0752),
				.a4(P0762),
				.a5(P0772),
				.a6(P0852),
				.a7(P0862),
				.a8(P0872),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02650)
);

assign C0650=c00650+c01650+c02650;
assign A0650=(C0650>=0)?1:0;

ninexnine_unit ninexnine_unit_270(
				.clk(clk),
				.rstn(rstn),
				.a0(P0660),
				.a1(P0670),
				.a2(P0680),
				.a3(P0760),
				.a4(P0770),
				.a5(P0780),
				.a6(P0860),
				.a7(P0870),
				.a8(P0880),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00660)
);

ninexnine_unit ninexnine_unit_271(
				.clk(clk),
				.rstn(rstn),
				.a0(P0661),
				.a1(P0671),
				.a2(P0681),
				.a3(P0761),
				.a4(P0771),
				.a5(P0781),
				.a6(P0861),
				.a7(P0871),
				.a8(P0881),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01660)
);

ninexnine_unit ninexnine_unit_272(
				.clk(clk),
				.rstn(rstn),
				.a0(P0662),
				.a1(P0672),
				.a2(P0682),
				.a3(P0762),
				.a4(P0772),
				.a5(P0782),
				.a6(P0862),
				.a7(P0872),
				.a8(P0882),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02660)
);

assign C0660=c00660+c01660+c02660;
assign A0660=(C0660>=0)?1:0;

ninexnine_unit ninexnine_unit_273(
				.clk(clk),
				.rstn(rstn),
				.a0(P0670),
				.a1(P0680),
				.a2(P0690),
				.a3(P0770),
				.a4(P0780),
				.a5(P0790),
				.a6(P0870),
				.a7(P0880),
				.a8(P0890),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00670)
);

ninexnine_unit ninexnine_unit_274(
				.clk(clk),
				.rstn(rstn),
				.a0(P0671),
				.a1(P0681),
				.a2(P0691),
				.a3(P0771),
				.a4(P0781),
				.a5(P0791),
				.a6(P0871),
				.a7(P0881),
				.a8(P0891),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01670)
);

ninexnine_unit ninexnine_unit_275(
				.clk(clk),
				.rstn(rstn),
				.a0(P0672),
				.a1(P0682),
				.a2(P0692),
				.a3(P0772),
				.a4(P0782),
				.a5(P0792),
				.a6(P0872),
				.a7(P0882),
				.a8(P0892),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02670)
);

assign C0670=c00670+c01670+c02670;
assign A0670=(C0670>=0)?1:0;

ninexnine_unit ninexnine_unit_276(
				.clk(clk),
				.rstn(rstn),
				.a0(P0680),
				.a1(P0690),
				.a2(P06A0),
				.a3(P0780),
				.a4(P0790),
				.a5(P07A0),
				.a6(P0880),
				.a7(P0890),
				.a8(P08A0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00680)
);

ninexnine_unit ninexnine_unit_277(
				.clk(clk),
				.rstn(rstn),
				.a0(P0681),
				.a1(P0691),
				.a2(P06A1),
				.a3(P0781),
				.a4(P0791),
				.a5(P07A1),
				.a6(P0881),
				.a7(P0891),
				.a8(P08A1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01680)
);

ninexnine_unit ninexnine_unit_278(
				.clk(clk),
				.rstn(rstn),
				.a0(P0682),
				.a1(P0692),
				.a2(P06A2),
				.a3(P0782),
				.a4(P0792),
				.a5(P07A2),
				.a6(P0882),
				.a7(P0892),
				.a8(P08A2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02680)
);

assign C0680=c00680+c01680+c02680;
assign A0680=(C0680>=0)?1:0;

ninexnine_unit ninexnine_unit_279(
				.clk(clk),
				.rstn(rstn),
				.a0(P0690),
				.a1(P06A0),
				.a2(P06B0),
				.a3(P0790),
				.a4(P07A0),
				.a5(P07B0),
				.a6(P0890),
				.a7(P08A0),
				.a8(P08B0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00690)
);

ninexnine_unit ninexnine_unit_280(
				.clk(clk),
				.rstn(rstn),
				.a0(P0691),
				.a1(P06A1),
				.a2(P06B1),
				.a3(P0791),
				.a4(P07A1),
				.a5(P07B1),
				.a6(P0891),
				.a7(P08A1),
				.a8(P08B1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01690)
);

ninexnine_unit ninexnine_unit_281(
				.clk(clk),
				.rstn(rstn),
				.a0(P0692),
				.a1(P06A2),
				.a2(P06B2),
				.a3(P0792),
				.a4(P07A2),
				.a5(P07B2),
				.a6(P0892),
				.a7(P08A2),
				.a8(P08B2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02690)
);

assign C0690=c00690+c01690+c02690;
assign A0690=(C0690>=0)?1:0;

ninexnine_unit ninexnine_unit_282(
				.clk(clk),
				.rstn(rstn),
				.a0(P06A0),
				.a1(P06B0),
				.a2(P06C0),
				.a3(P07A0),
				.a4(P07B0),
				.a5(P07C0),
				.a6(P08A0),
				.a7(P08B0),
				.a8(P08C0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c006A0)
);

ninexnine_unit ninexnine_unit_283(
				.clk(clk),
				.rstn(rstn),
				.a0(P06A1),
				.a1(P06B1),
				.a2(P06C1),
				.a3(P07A1),
				.a4(P07B1),
				.a5(P07C1),
				.a6(P08A1),
				.a7(P08B1),
				.a8(P08C1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c016A0)
);

ninexnine_unit ninexnine_unit_284(
				.clk(clk),
				.rstn(rstn),
				.a0(P06A2),
				.a1(P06B2),
				.a2(P06C2),
				.a3(P07A2),
				.a4(P07B2),
				.a5(P07C2),
				.a6(P08A2),
				.a7(P08B2),
				.a8(P08C2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c026A0)
);

assign C06A0=c006A0+c016A0+c026A0;
assign A06A0=(C06A0>=0)?1:0;

ninexnine_unit ninexnine_unit_285(
				.clk(clk),
				.rstn(rstn),
				.a0(P06B0),
				.a1(P06C0),
				.a2(P06D0),
				.a3(P07B0),
				.a4(P07C0),
				.a5(P07D0),
				.a6(P08B0),
				.a7(P08C0),
				.a8(P08D0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c006B0)
);

ninexnine_unit ninexnine_unit_286(
				.clk(clk),
				.rstn(rstn),
				.a0(P06B1),
				.a1(P06C1),
				.a2(P06D1),
				.a3(P07B1),
				.a4(P07C1),
				.a5(P07D1),
				.a6(P08B1),
				.a7(P08C1),
				.a8(P08D1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c016B0)
);

ninexnine_unit ninexnine_unit_287(
				.clk(clk),
				.rstn(rstn),
				.a0(P06B2),
				.a1(P06C2),
				.a2(P06D2),
				.a3(P07B2),
				.a4(P07C2),
				.a5(P07D2),
				.a6(P08B2),
				.a7(P08C2),
				.a8(P08D2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c026B0)
);

assign C06B0=c006B0+c016B0+c026B0;
assign A06B0=(C06B0>=0)?1:0;

ninexnine_unit ninexnine_unit_288(
				.clk(clk),
				.rstn(rstn),
				.a0(P06C0),
				.a1(P06D0),
				.a2(P06E0),
				.a3(P07C0),
				.a4(P07D0),
				.a5(P07E0),
				.a6(P08C0),
				.a7(P08D0),
				.a8(P08E0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c006C0)
);

ninexnine_unit ninexnine_unit_289(
				.clk(clk),
				.rstn(rstn),
				.a0(P06C1),
				.a1(P06D1),
				.a2(P06E1),
				.a3(P07C1),
				.a4(P07D1),
				.a5(P07E1),
				.a6(P08C1),
				.a7(P08D1),
				.a8(P08E1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c016C0)
);

ninexnine_unit ninexnine_unit_290(
				.clk(clk),
				.rstn(rstn),
				.a0(P06C2),
				.a1(P06D2),
				.a2(P06E2),
				.a3(P07C2),
				.a4(P07D2),
				.a5(P07E2),
				.a6(P08C2),
				.a7(P08D2),
				.a8(P08E2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c026C0)
);

assign C06C0=c006C0+c016C0+c026C0;
assign A06C0=(C06C0>=0)?1:0;

ninexnine_unit ninexnine_unit_291(
				.clk(clk),
				.rstn(rstn),
				.a0(P06D0),
				.a1(P06E0),
				.a2(P06F0),
				.a3(P07D0),
				.a4(P07E0),
				.a5(P07F0),
				.a6(P08D0),
				.a7(P08E0),
				.a8(P08F0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c006D0)
);

ninexnine_unit ninexnine_unit_292(
				.clk(clk),
				.rstn(rstn),
				.a0(P06D1),
				.a1(P06E1),
				.a2(P06F1),
				.a3(P07D1),
				.a4(P07E1),
				.a5(P07F1),
				.a6(P08D1),
				.a7(P08E1),
				.a8(P08F1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c016D0)
);

ninexnine_unit ninexnine_unit_293(
				.clk(clk),
				.rstn(rstn),
				.a0(P06D2),
				.a1(P06E2),
				.a2(P06F2),
				.a3(P07D2),
				.a4(P07E2),
				.a5(P07F2),
				.a6(P08D2),
				.a7(P08E2),
				.a8(P08F2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c026D0)
);

assign C06D0=c006D0+c016D0+c026D0;
assign A06D0=(C06D0>=0)?1:0;

ninexnine_unit ninexnine_unit_294(
				.clk(clk),
				.rstn(rstn),
				.a0(P0700),
				.a1(P0710),
				.a2(P0720),
				.a3(P0800),
				.a4(P0810),
				.a5(P0820),
				.a6(P0900),
				.a7(P0910),
				.a8(P0920),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00700)
);

ninexnine_unit ninexnine_unit_295(
				.clk(clk),
				.rstn(rstn),
				.a0(P0701),
				.a1(P0711),
				.a2(P0721),
				.a3(P0801),
				.a4(P0811),
				.a5(P0821),
				.a6(P0901),
				.a7(P0911),
				.a8(P0921),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01700)
);

ninexnine_unit ninexnine_unit_296(
				.clk(clk),
				.rstn(rstn),
				.a0(P0702),
				.a1(P0712),
				.a2(P0722),
				.a3(P0802),
				.a4(P0812),
				.a5(P0822),
				.a6(P0902),
				.a7(P0912),
				.a8(P0922),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02700)
);

assign C0700=c00700+c01700+c02700;
assign A0700=(C0700>=0)?1:0;

ninexnine_unit ninexnine_unit_297(
				.clk(clk),
				.rstn(rstn),
				.a0(P0710),
				.a1(P0720),
				.a2(P0730),
				.a3(P0810),
				.a4(P0820),
				.a5(P0830),
				.a6(P0910),
				.a7(P0920),
				.a8(P0930),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00710)
);

ninexnine_unit ninexnine_unit_298(
				.clk(clk),
				.rstn(rstn),
				.a0(P0711),
				.a1(P0721),
				.a2(P0731),
				.a3(P0811),
				.a4(P0821),
				.a5(P0831),
				.a6(P0911),
				.a7(P0921),
				.a8(P0931),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01710)
);

ninexnine_unit ninexnine_unit_299(
				.clk(clk),
				.rstn(rstn),
				.a0(P0712),
				.a1(P0722),
				.a2(P0732),
				.a3(P0812),
				.a4(P0822),
				.a5(P0832),
				.a6(P0912),
				.a7(P0922),
				.a8(P0932),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02710)
);

assign C0710=c00710+c01710+c02710;
assign A0710=(C0710>=0)?1:0;

ninexnine_unit ninexnine_unit_300(
				.clk(clk),
				.rstn(rstn),
				.a0(P0720),
				.a1(P0730),
				.a2(P0740),
				.a3(P0820),
				.a4(P0830),
				.a5(P0840),
				.a6(P0920),
				.a7(P0930),
				.a8(P0940),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00720)
);

ninexnine_unit ninexnine_unit_301(
				.clk(clk),
				.rstn(rstn),
				.a0(P0721),
				.a1(P0731),
				.a2(P0741),
				.a3(P0821),
				.a4(P0831),
				.a5(P0841),
				.a6(P0921),
				.a7(P0931),
				.a8(P0941),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01720)
);

ninexnine_unit ninexnine_unit_302(
				.clk(clk),
				.rstn(rstn),
				.a0(P0722),
				.a1(P0732),
				.a2(P0742),
				.a3(P0822),
				.a4(P0832),
				.a5(P0842),
				.a6(P0922),
				.a7(P0932),
				.a8(P0942),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02720)
);

assign C0720=c00720+c01720+c02720;
assign A0720=(C0720>=0)?1:0;

ninexnine_unit ninexnine_unit_303(
				.clk(clk),
				.rstn(rstn),
				.a0(P0730),
				.a1(P0740),
				.a2(P0750),
				.a3(P0830),
				.a4(P0840),
				.a5(P0850),
				.a6(P0930),
				.a7(P0940),
				.a8(P0950),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00730)
);

ninexnine_unit ninexnine_unit_304(
				.clk(clk),
				.rstn(rstn),
				.a0(P0731),
				.a1(P0741),
				.a2(P0751),
				.a3(P0831),
				.a4(P0841),
				.a5(P0851),
				.a6(P0931),
				.a7(P0941),
				.a8(P0951),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01730)
);

ninexnine_unit ninexnine_unit_305(
				.clk(clk),
				.rstn(rstn),
				.a0(P0732),
				.a1(P0742),
				.a2(P0752),
				.a3(P0832),
				.a4(P0842),
				.a5(P0852),
				.a6(P0932),
				.a7(P0942),
				.a8(P0952),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02730)
);

assign C0730=c00730+c01730+c02730;
assign A0730=(C0730>=0)?1:0;

ninexnine_unit ninexnine_unit_306(
				.clk(clk),
				.rstn(rstn),
				.a0(P0740),
				.a1(P0750),
				.a2(P0760),
				.a3(P0840),
				.a4(P0850),
				.a5(P0860),
				.a6(P0940),
				.a7(P0950),
				.a8(P0960),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00740)
);

ninexnine_unit ninexnine_unit_307(
				.clk(clk),
				.rstn(rstn),
				.a0(P0741),
				.a1(P0751),
				.a2(P0761),
				.a3(P0841),
				.a4(P0851),
				.a5(P0861),
				.a6(P0941),
				.a7(P0951),
				.a8(P0961),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01740)
);

ninexnine_unit ninexnine_unit_308(
				.clk(clk),
				.rstn(rstn),
				.a0(P0742),
				.a1(P0752),
				.a2(P0762),
				.a3(P0842),
				.a4(P0852),
				.a5(P0862),
				.a6(P0942),
				.a7(P0952),
				.a8(P0962),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02740)
);

assign C0740=c00740+c01740+c02740;
assign A0740=(C0740>=0)?1:0;

ninexnine_unit ninexnine_unit_309(
				.clk(clk),
				.rstn(rstn),
				.a0(P0750),
				.a1(P0760),
				.a2(P0770),
				.a3(P0850),
				.a4(P0860),
				.a5(P0870),
				.a6(P0950),
				.a7(P0960),
				.a8(P0970),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00750)
);

ninexnine_unit ninexnine_unit_310(
				.clk(clk),
				.rstn(rstn),
				.a0(P0751),
				.a1(P0761),
				.a2(P0771),
				.a3(P0851),
				.a4(P0861),
				.a5(P0871),
				.a6(P0951),
				.a7(P0961),
				.a8(P0971),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01750)
);

ninexnine_unit ninexnine_unit_311(
				.clk(clk),
				.rstn(rstn),
				.a0(P0752),
				.a1(P0762),
				.a2(P0772),
				.a3(P0852),
				.a4(P0862),
				.a5(P0872),
				.a6(P0952),
				.a7(P0962),
				.a8(P0972),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02750)
);

assign C0750=c00750+c01750+c02750;
assign A0750=(C0750>=0)?1:0;

ninexnine_unit ninexnine_unit_312(
				.clk(clk),
				.rstn(rstn),
				.a0(P0760),
				.a1(P0770),
				.a2(P0780),
				.a3(P0860),
				.a4(P0870),
				.a5(P0880),
				.a6(P0960),
				.a7(P0970),
				.a8(P0980),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00760)
);

ninexnine_unit ninexnine_unit_313(
				.clk(clk),
				.rstn(rstn),
				.a0(P0761),
				.a1(P0771),
				.a2(P0781),
				.a3(P0861),
				.a4(P0871),
				.a5(P0881),
				.a6(P0961),
				.a7(P0971),
				.a8(P0981),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01760)
);

ninexnine_unit ninexnine_unit_314(
				.clk(clk),
				.rstn(rstn),
				.a0(P0762),
				.a1(P0772),
				.a2(P0782),
				.a3(P0862),
				.a4(P0872),
				.a5(P0882),
				.a6(P0962),
				.a7(P0972),
				.a8(P0982),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02760)
);

assign C0760=c00760+c01760+c02760;
assign A0760=(C0760>=0)?1:0;

ninexnine_unit ninexnine_unit_315(
				.clk(clk),
				.rstn(rstn),
				.a0(P0770),
				.a1(P0780),
				.a2(P0790),
				.a3(P0870),
				.a4(P0880),
				.a5(P0890),
				.a6(P0970),
				.a7(P0980),
				.a8(P0990),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00770)
);

ninexnine_unit ninexnine_unit_316(
				.clk(clk),
				.rstn(rstn),
				.a0(P0771),
				.a1(P0781),
				.a2(P0791),
				.a3(P0871),
				.a4(P0881),
				.a5(P0891),
				.a6(P0971),
				.a7(P0981),
				.a8(P0991),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01770)
);

ninexnine_unit ninexnine_unit_317(
				.clk(clk),
				.rstn(rstn),
				.a0(P0772),
				.a1(P0782),
				.a2(P0792),
				.a3(P0872),
				.a4(P0882),
				.a5(P0892),
				.a6(P0972),
				.a7(P0982),
				.a8(P0992),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02770)
);

assign C0770=c00770+c01770+c02770;
assign A0770=(C0770>=0)?1:0;

ninexnine_unit ninexnine_unit_318(
				.clk(clk),
				.rstn(rstn),
				.a0(P0780),
				.a1(P0790),
				.a2(P07A0),
				.a3(P0880),
				.a4(P0890),
				.a5(P08A0),
				.a6(P0980),
				.a7(P0990),
				.a8(P09A0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00780)
);

ninexnine_unit ninexnine_unit_319(
				.clk(clk),
				.rstn(rstn),
				.a0(P0781),
				.a1(P0791),
				.a2(P07A1),
				.a3(P0881),
				.a4(P0891),
				.a5(P08A1),
				.a6(P0981),
				.a7(P0991),
				.a8(P09A1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01780)
);

ninexnine_unit ninexnine_unit_320(
				.clk(clk),
				.rstn(rstn),
				.a0(P0782),
				.a1(P0792),
				.a2(P07A2),
				.a3(P0882),
				.a4(P0892),
				.a5(P08A2),
				.a6(P0982),
				.a7(P0992),
				.a8(P09A2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02780)
);

assign C0780=c00780+c01780+c02780;
assign A0780=(C0780>=0)?1:0;

ninexnine_unit ninexnine_unit_321(
				.clk(clk),
				.rstn(rstn),
				.a0(P0790),
				.a1(P07A0),
				.a2(P07B0),
				.a3(P0890),
				.a4(P08A0),
				.a5(P08B0),
				.a6(P0990),
				.a7(P09A0),
				.a8(P09B0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00790)
);

ninexnine_unit ninexnine_unit_322(
				.clk(clk),
				.rstn(rstn),
				.a0(P0791),
				.a1(P07A1),
				.a2(P07B1),
				.a3(P0891),
				.a4(P08A1),
				.a5(P08B1),
				.a6(P0991),
				.a7(P09A1),
				.a8(P09B1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01790)
);

ninexnine_unit ninexnine_unit_323(
				.clk(clk),
				.rstn(rstn),
				.a0(P0792),
				.a1(P07A2),
				.a2(P07B2),
				.a3(P0892),
				.a4(P08A2),
				.a5(P08B2),
				.a6(P0992),
				.a7(P09A2),
				.a8(P09B2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02790)
);

assign C0790=c00790+c01790+c02790;
assign A0790=(C0790>=0)?1:0;

ninexnine_unit ninexnine_unit_324(
				.clk(clk),
				.rstn(rstn),
				.a0(P07A0),
				.a1(P07B0),
				.a2(P07C0),
				.a3(P08A0),
				.a4(P08B0),
				.a5(P08C0),
				.a6(P09A0),
				.a7(P09B0),
				.a8(P09C0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c007A0)
);

ninexnine_unit ninexnine_unit_325(
				.clk(clk),
				.rstn(rstn),
				.a0(P07A1),
				.a1(P07B1),
				.a2(P07C1),
				.a3(P08A1),
				.a4(P08B1),
				.a5(P08C1),
				.a6(P09A1),
				.a7(P09B1),
				.a8(P09C1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c017A0)
);

ninexnine_unit ninexnine_unit_326(
				.clk(clk),
				.rstn(rstn),
				.a0(P07A2),
				.a1(P07B2),
				.a2(P07C2),
				.a3(P08A2),
				.a4(P08B2),
				.a5(P08C2),
				.a6(P09A2),
				.a7(P09B2),
				.a8(P09C2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c027A0)
);

assign C07A0=c007A0+c017A0+c027A0;
assign A07A0=(C07A0>=0)?1:0;

ninexnine_unit ninexnine_unit_327(
				.clk(clk),
				.rstn(rstn),
				.a0(P07B0),
				.a1(P07C0),
				.a2(P07D0),
				.a3(P08B0),
				.a4(P08C0),
				.a5(P08D0),
				.a6(P09B0),
				.a7(P09C0),
				.a8(P09D0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c007B0)
);

ninexnine_unit ninexnine_unit_328(
				.clk(clk),
				.rstn(rstn),
				.a0(P07B1),
				.a1(P07C1),
				.a2(P07D1),
				.a3(P08B1),
				.a4(P08C1),
				.a5(P08D1),
				.a6(P09B1),
				.a7(P09C1),
				.a8(P09D1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c017B0)
);

ninexnine_unit ninexnine_unit_329(
				.clk(clk),
				.rstn(rstn),
				.a0(P07B2),
				.a1(P07C2),
				.a2(P07D2),
				.a3(P08B2),
				.a4(P08C2),
				.a5(P08D2),
				.a6(P09B2),
				.a7(P09C2),
				.a8(P09D2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c027B0)
);

assign C07B0=c007B0+c017B0+c027B0;
assign A07B0=(C07B0>=0)?1:0;

ninexnine_unit ninexnine_unit_330(
				.clk(clk),
				.rstn(rstn),
				.a0(P07C0),
				.a1(P07D0),
				.a2(P07E0),
				.a3(P08C0),
				.a4(P08D0),
				.a5(P08E0),
				.a6(P09C0),
				.a7(P09D0),
				.a8(P09E0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c007C0)
);

ninexnine_unit ninexnine_unit_331(
				.clk(clk),
				.rstn(rstn),
				.a0(P07C1),
				.a1(P07D1),
				.a2(P07E1),
				.a3(P08C1),
				.a4(P08D1),
				.a5(P08E1),
				.a6(P09C1),
				.a7(P09D1),
				.a8(P09E1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c017C0)
);

ninexnine_unit ninexnine_unit_332(
				.clk(clk),
				.rstn(rstn),
				.a0(P07C2),
				.a1(P07D2),
				.a2(P07E2),
				.a3(P08C2),
				.a4(P08D2),
				.a5(P08E2),
				.a6(P09C2),
				.a7(P09D2),
				.a8(P09E2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c027C0)
);

assign C07C0=c007C0+c017C0+c027C0;
assign A07C0=(C07C0>=0)?1:0;

ninexnine_unit ninexnine_unit_333(
				.clk(clk),
				.rstn(rstn),
				.a0(P07D0),
				.a1(P07E0),
				.a2(P07F0),
				.a3(P08D0),
				.a4(P08E0),
				.a5(P08F0),
				.a6(P09D0),
				.a7(P09E0),
				.a8(P09F0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c007D0)
);

ninexnine_unit ninexnine_unit_334(
				.clk(clk),
				.rstn(rstn),
				.a0(P07D1),
				.a1(P07E1),
				.a2(P07F1),
				.a3(P08D1),
				.a4(P08E1),
				.a5(P08F1),
				.a6(P09D1),
				.a7(P09E1),
				.a8(P09F1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c017D0)
);

ninexnine_unit ninexnine_unit_335(
				.clk(clk),
				.rstn(rstn),
				.a0(P07D2),
				.a1(P07E2),
				.a2(P07F2),
				.a3(P08D2),
				.a4(P08E2),
				.a5(P08F2),
				.a6(P09D2),
				.a7(P09E2),
				.a8(P09F2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c027D0)
);

assign C07D0=c007D0+c017D0+c027D0;
assign A07D0=(C07D0>=0)?1:0;

ninexnine_unit ninexnine_unit_336(
				.clk(clk),
				.rstn(rstn),
				.a0(P0800),
				.a1(P0810),
				.a2(P0820),
				.a3(P0900),
				.a4(P0910),
				.a5(P0920),
				.a6(P0A00),
				.a7(P0A10),
				.a8(P0A20),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00800)
);

ninexnine_unit ninexnine_unit_337(
				.clk(clk),
				.rstn(rstn),
				.a0(P0801),
				.a1(P0811),
				.a2(P0821),
				.a3(P0901),
				.a4(P0911),
				.a5(P0921),
				.a6(P0A01),
				.a7(P0A11),
				.a8(P0A21),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01800)
);

ninexnine_unit ninexnine_unit_338(
				.clk(clk),
				.rstn(rstn),
				.a0(P0802),
				.a1(P0812),
				.a2(P0822),
				.a3(P0902),
				.a4(P0912),
				.a5(P0922),
				.a6(P0A02),
				.a7(P0A12),
				.a8(P0A22),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02800)
);

assign C0800=c00800+c01800+c02800;
assign A0800=(C0800>=0)?1:0;

ninexnine_unit ninexnine_unit_339(
				.clk(clk),
				.rstn(rstn),
				.a0(P0810),
				.a1(P0820),
				.a2(P0830),
				.a3(P0910),
				.a4(P0920),
				.a5(P0930),
				.a6(P0A10),
				.a7(P0A20),
				.a8(P0A30),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00810)
);

ninexnine_unit ninexnine_unit_340(
				.clk(clk),
				.rstn(rstn),
				.a0(P0811),
				.a1(P0821),
				.a2(P0831),
				.a3(P0911),
				.a4(P0921),
				.a5(P0931),
				.a6(P0A11),
				.a7(P0A21),
				.a8(P0A31),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01810)
);

ninexnine_unit ninexnine_unit_341(
				.clk(clk),
				.rstn(rstn),
				.a0(P0812),
				.a1(P0822),
				.a2(P0832),
				.a3(P0912),
				.a4(P0922),
				.a5(P0932),
				.a6(P0A12),
				.a7(P0A22),
				.a8(P0A32),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02810)
);

assign C0810=c00810+c01810+c02810;
assign A0810=(C0810>=0)?1:0;

ninexnine_unit ninexnine_unit_342(
				.clk(clk),
				.rstn(rstn),
				.a0(P0820),
				.a1(P0830),
				.a2(P0840),
				.a3(P0920),
				.a4(P0930),
				.a5(P0940),
				.a6(P0A20),
				.a7(P0A30),
				.a8(P0A40),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00820)
);

ninexnine_unit ninexnine_unit_343(
				.clk(clk),
				.rstn(rstn),
				.a0(P0821),
				.a1(P0831),
				.a2(P0841),
				.a3(P0921),
				.a4(P0931),
				.a5(P0941),
				.a6(P0A21),
				.a7(P0A31),
				.a8(P0A41),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01820)
);

ninexnine_unit ninexnine_unit_344(
				.clk(clk),
				.rstn(rstn),
				.a0(P0822),
				.a1(P0832),
				.a2(P0842),
				.a3(P0922),
				.a4(P0932),
				.a5(P0942),
				.a6(P0A22),
				.a7(P0A32),
				.a8(P0A42),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02820)
);

assign C0820=c00820+c01820+c02820;
assign A0820=(C0820>=0)?1:0;

ninexnine_unit ninexnine_unit_345(
				.clk(clk),
				.rstn(rstn),
				.a0(P0830),
				.a1(P0840),
				.a2(P0850),
				.a3(P0930),
				.a4(P0940),
				.a5(P0950),
				.a6(P0A30),
				.a7(P0A40),
				.a8(P0A50),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00830)
);

ninexnine_unit ninexnine_unit_346(
				.clk(clk),
				.rstn(rstn),
				.a0(P0831),
				.a1(P0841),
				.a2(P0851),
				.a3(P0931),
				.a4(P0941),
				.a5(P0951),
				.a6(P0A31),
				.a7(P0A41),
				.a8(P0A51),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01830)
);

ninexnine_unit ninexnine_unit_347(
				.clk(clk),
				.rstn(rstn),
				.a0(P0832),
				.a1(P0842),
				.a2(P0852),
				.a3(P0932),
				.a4(P0942),
				.a5(P0952),
				.a6(P0A32),
				.a7(P0A42),
				.a8(P0A52),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02830)
);

assign C0830=c00830+c01830+c02830;
assign A0830=(C0830>=0)?1:0;

ninexnine_unit ninexnine_unit_348(
				.clk(clk),
				.rstn(rstn),
				.a0(P0840),
				.a1(P0850),
				.a2(P0860),
				.a3(P0940),
				.a4(P0950),
				.a5(P0960),
				.a6(P0A40),
				.a7(P0A50),
				.a8(P0A60),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00840)
);

ninexnine_unit ninexnine_unit_349(
				.clk(clk),
				.rstn(rstn),
				.a0(P0841),
				.a1(P0851),
				.a2(P0861),
				.a3(P0941),
				.a4(P0951),
				.a5(P0961),
				.a6(P0A41),
				.a7(P0A51),
				.a8(P0A61),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01840)
);

ninexnine_unit ninexnine_unit_350(
				.clk(clk),
				.rstn(rstn),
				.a0(P0842),
				.a1(P0852),
				.a2(P0862),
				.a3(P0942),
				.a4(P0952),
				.a5(P0962),
				.a6(P0A42),
				.a7(P0A52),
				.a8(P0A62),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02840)
);

assign C0840=c00840+c01840+c02840;
assign A0840=(C0840>=0)?1:0;

ninexnine_unit ninexnine_unit_351(
				.clk(clk),
				.rstn(rstn),
				.a0(P0850),
				.a1(P0860),
				.a2(P0870),
				.a3(P0950),
				.a4(P0960),
				.a5(P0970),
				.a6(P0A50),
				.a7(P0A60),
				.a8(P0A70),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00850)
);

ninexnine_unit ninexnine_unit_352(
				.clk(clk),
				.rstn(rstn),
				.a0(P0851),
				.a1(P0861),
				.a2(P0871),
				.a3(P0951),
				.a4(P0961),
				.a5(P0971),
				.a6(P0A51),
				.a7(P0A61),
				.a8(P0A71),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01850)
);

ninexnine_unit ninexnine_unit_353(
				.clk(clk),
				.rstn(rstn),
				.a0(P0852),
				.a1(P0862),
				.a2(P0872),
				.a3(P0952),
				.a4(P0962),
				.a5(P0972),
				.a6(P0A52),
				.a7(P0A62),
				.a8(P0A72),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02850)
);

assign C0850=c00850+c01850+c02850;
assign A0850=(C0850>=0)?1:0;

ninexnine_unit ninexnine_unit_354(
				.clk(clk),
				.rstn(rstn),
				.a0(P0860),
				.a1(P0870),
				.a2(P0880),
				.a3(P0960),
				.a4(P0970),
				.a5(P0980),
				.a6(P0A60),
				.a7(P0A70),
				.a8(P0A80),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00860)
);

ninexnine_unit ninexnine_unit_355(
				.clk(clk),
				.rstn(rstn),
				.a0(P0861),
				.a1(P0871),
				.a2(P0881),
				.a3(P0961),
				.a4(P0971),
				.a5(P0981),
				.a6(P0A61),
				.a7(P0A71),
				.a8(P0A81),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01860)
);

ninexnine_unit ninexnine_unit_356(
				.clk(clk),
				.rstn(rstn),
				.a0(P0862),
				.a1(P0872),
				.a2(P0882),
				.a3(P0962),
				.a4(P0972),
				.a5(P0982),
				.a6(P0A62),
				.a7(P0A72),
				.a8(P0A82),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02860)
);

assign C0860=c00860+c01860+c02860;
assign A0860=(C0860>=0)?1:0;

ninexnine_unit ninexnine_unit_357(
				.clk(clk),
				.rstn(rstn),
				.a0(P0870),
				.a1(P0880),
				.a2(P0890),
				.a3(P0970),
				.a4(P0980),
				.a5(P0990),
				.a6(P0A70),
				.a7(P0A80),
				.a8(P0A90),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00870)
);

ninexnine_unit ninexnine_unit_358(
				.clk(clk),
				.rstn(rstn),
				.a0(P0871),
				.a1(P0881),
				.a2(P0891),
				.a3(P0971),
				.a4(P0981),
				.a5(P0991),
				.a6(P0A71),
				.a7(P0A81),
				.a8(P0A91),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01870)
);

ninexnine_unit ninexnine_unit_359(
				.clk(clk),
				.rstn(rstn),
				.a0(P0872),
				.a1(P0882),
				.a2(P0892),
				.a3(P0972),
				.a4(P0982),
				.a5(P0992),
				.a6(P0A72),
				.a7(P0A82),
				.a8(P0A92),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02870)
);

assign C0870=c00870+c01870+c02870;
assign A0870=(C0870>=0)?1:0;

ninexnine_unit ninexnine_unit_360(
				.clk(clk),
				.rstn(rstn),
				.a0(P0880),
				.a1(P0890),
				.a2(P08A0),
				.a3(P0980),
				.a4(P0990),
				.a5(P09A0),
				.a6(P0A80),
				.a7(P0A90),
				.a8(P0AA0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00880)
);

ninexnine_unit ninexnine_unit_361(
				.clk(clk),
				.rstn(rstn),
				.a0(P0881),
				.a1(P0891),
				.a2(P08A1),
				.a3(P0981),
				.a4(P0991),
				.a5(P09A1),
				.a6(P0A81),
				.a7(P0A91),
				.a8(P0AA1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01880)
);

ninexnine_unit ninexnine_unit_362(
				.clk(clk),
				.rstn(rstn),
				.a0(P0882),
				.a1(P0892),
				.a2(P08A2),
				.a3(P0982),
				.a4(P0992),
				.a5(P09A2),
				.a6(P0A82),
				.a7(P0A92),
				.a8(P0AA2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02880)
);

assign C0880=c00880+c01880+c02880;
assign A0880=(C0880>=0)?1:0;

ninexnine_unit ninexnine_unit_363(
				.clk(clk),
				.rstn(rstn),
				.a0(P0890),
				.a1(P08A0),
				.a2(P08B0),
				.a3(P0990),
				.a4(P09A0),
				.a5(P09B0),
				.a6(P0A90),
				.a7(P0AA0),
				.a8(P0AB0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00890)
);

ninexnine_unit ninexnine_unit_364(
				.clk(clk),
				.rstn(rstn),
				.a0(P0891),
				.a1(P08A1),
				.a2(P08B1),
				.a3(P0991),
				.a4(P09A1),
				.a5(P09B1),
				.a6(P0A91),
				.a7(P0AA1),
				.a8(P0AB1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01890)
);

ninexnine_unit ninexnine_unit_365(
				.clk(clk),
				.rstn(rstn),
				.a0(P0892),
				.a1(P08A2),
				.a2(P08B2),
				.a3(P0992),
				.a4(P09A2),
				.a5(P09B2),
				.a6(P0A92),
				.a7(P0AA2),
				.a8(P0AB2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02890)
);

assign C0890=c00890+c01890+c02890;
assign A0890=(C0890>=0)?1:0;

ninexnine_unit ninexnine_unit_366(
				.clk(clk),
				.rstn(rstn),
				.a0(P08A0),
				.a1(P08B0),
				.a2(P08C0),
				.a3(P09A0),
				.a4(P09B0),
				.a5(P09C0),
				.a6(P0AA0),
				.a7(P0AB0),
				.a8(P0AC0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c008A0)
);

ninexnine_unit ninexnine_unit_367(
				.clk(clk),
				.rstn(rstn),
				.a0(P08A1),
				.a1(P08B1),
				.a2(P08C1),
				.a3(P09A1),
				.a4(P09B1),
				.a5(P09C1),
				.a6(P0AA1),
				.a7(P0AB1),
				.a8(P0AC1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c018A0)
);

ninexnine_unit ninexnine_unit_368(
				.clk(clk),
				.rstn(rstn),
				.a0(P08A2),
				.a1(P08B2),
				.a2(P08C2),
				.a3(P09A2),
				.a4(P09B2),
				.a5(P09C2),
				.a6(P0AA2),
				.a7(P0AB2),
				.a8(P0AC2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c028A0)
);

assign C08A0=c008A0+c018A0+c028A0;
assign A08A0=(C08A0>=0)?1:0;

ninexnine_unit ninexnine_unit_369(
				.clk(clk),
				.rstn(rstn),
				.a0(P08B0),
				.a1(P08C0),
				.a2(P08D0),
				.a3(P09B0),
				.a4(P09C0),
				.a5(P09D0),
				.a6(P0AB0),
				.a7(P0AC0),
				.a8(P0AD0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c008B0)
);

ninexnine_unit ninexnine_unit_370(
				.clk(clk),
				.rstn(rstn),
				.a0(P08B1),
				.a1(P08C1),
				.a2(P08D1),
				.a3(P09B1),
				.a4(P09C1),
				.a5(P09D1),
				.a6(P0AB1),
				.a7(P0AC1),
				.a8(P0AD1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c018B0)
);

ninexnine_unit ninexnine_unit_371(
				.clk(clk),
				.rstn(rstn),
				.a0(P08B2),
				.a1(P08C2),
				.a2(P08D2),
				.a3(P09B2),
				.a4(P09C2),
				.a5(P09D2),
				.a6(P0AB2),
				.a7(P0AC2),
				.a8(P0AD2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c028B0)
);

assign C08B0=c008B0+c018B0+c028B0;
assign A08B0=(C08B0>=0)?1:0;

ninexnine_unit ninexnine_unit_372(
				.clk(clk),
				.rstn(rstn),
				.a0(P08C0),
				.a1(P08D0),
				.a2(P08E0),
				.a3(P09C0),
				.a4(P09D0),
				.a5(P09E0),
				.a6(P0AC0),
				.a7(P0AD0),
				.a8(P0AE0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c008C0)
);

ninexnine_unit ninexnine_unit_373(
				.clk(clk),
				.rstn(rstn),
				.a0(P08C1),
				.a1(P08D1),
				.a2(P08E1),
				.a3(P09C1),
				.a4(P09D1),
				.a5(P09E1),
				.a6(P0AC1),
				.a7(P0AD1),
				.a8(P0AE1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c018C0)
);

ninexnine_unit ninexnine_unit_374(
				.clk(clk),
				.rstn(rstn),
				.a0(P08C2),
				.a1(P08D2),
				.a2(P08E2),
				.a3(P09C2),
				.a4(P09D2),
				.a5(P09E2),
				.a6(P0AC2),
				.a7(P0AD2),
				.a8(P0AE2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c028C0)
);

assign C08C0=c008C0+c018C0+c028C0;
assign A08C0=(C08C0>=0)?1:0;

ninexnine_unit ninexnine_unit_375(
				.clk(clk),
				.rstn(rstn),
				.a0(P08D0),
				.a1(P08E0),
				.a2(P08F0),
				.a3(P09D0),
				.a4(P09E0),
				.a5(P09F0),
				.a6(P0AD0),
				.a7(P0AE0),
				.a8(P0AF0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c008D0)
);

ninexnine_unit ninexnine_unit_376(
				.clk(clk),
				.rstn(rstn),
				.a0(P08D1),
				.a1(P08E1),
				.a2(P08F1),
				.a3(P09D1),
				.a4(P09E1),
				.a5(P09F1),
				.a6(P0AD1),
				.a7(P0AE1),
				.a8(P0AF1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c018D0)
);

ninexnine_unit ninexnine_unit_377(
				.clk(clk),
				.rstn(rstn),
				.a0(P08D2),
				.a1(P08E2),
				.a2(P08F2),
				.a3(P09D2),
				.a4(P09E2),
				.a5(P09F2),
				.a6(P0AD2),
				.a7(P0AE2),
				.a8(P0AF2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c028D0)
);

assign C08D0=c008D0+c018D0+c028D0;
assign A08D0=(C08D0>=0)?1:0;

ninexnine_unit ninexnine_unit_378(
				.clk(clk),
				.rstn(rstn),
				.a0(P0900),
				.a1(P0910),
				.a2(P0920),
				.a3(P0A00),
				.a4(P0A10),
				.a5(P0A20),
				.a6(P0B00),
				.a7(P0B10),
				.a8(P0B20),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00900)
);

ninexnine_unit ninexnine_unit_379(
				.clk(clk),
				.rstn(rstn),
				.a0(P0901),
				.a1(P0911),
				.a2(P0921),
				.a3(P0A01),
				.a4(P0A11),
				.a5(P0A21),
				.a6(P0B01),
				.a7(P0B11),
				.a8(P0B21),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01900)
);

ninexnine_unit ninexnine_unit_380(
				.clk(clk),
				.rstn(rstn),
				.a0(P0902),
				.a1(P0912),
				.a2(P0922),
				.a3(P0A02),
				.a4(P0A12),
				.a5(P0A22),
				.a6(P0B02),
				.a7(P0B12),
				.a8(P0B22),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02900)
);

assign C0900=c00900+c01900+c02900;
assign A0900=(C0900>=0)?1:0;

ninexnine_unit ninexnine_unit_381(
				.clk(clk),
				.rstn(rstn),
				.a0(P0910),
				.a1(P0920),
				.a2(P0930),
				.a3(P0A10),
				.a4(P0A20),
				.a5(P0A30),
				.a6(P0B10),
				.a7(P0B20),
				.a8(P0B30),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00910)
);

ninexnine_unit ninexnine_unit_382(
				.clk(clk),
				.rstn(rstn),
				.a0(P0911),
				.a1(P0921),
				.a2(P0931),
				.a3(P0A11),
				.a4(P0A21),
				.a5(P0A31),
				.a6(P0B11),
				.a7(P0B21),
				.a8(P0B31),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01910)
);

ninexnine_unit ninexnine_unit_383(
				.clk(clk),
				.rstn(rstn),
				.a0(P0912),
				.a1(P0922),
				.a2(P0932),
				.a3(P0A12),
				.a4(P0A22),
				.a5(P0A32),
				.a6(P0B12),
				.a7(P0B22),
				.a8(P0B32),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02910)
);

assign C0910=c00910+c01910+c02910;
assign A0910=(C0910>=0)?1:0;

ninexnine_unit ninexnine_unit_384(
				.clk(clk),
				.rstn(rstn),
				.a0(P0920),
				.a1(P0930),
				.a2(P0940),
				.a3(P0A20),
				.a4(P0A30),
				.a5(P0A40),
				.a6(P0B20),
				.a7(P0B30),
				.a8(P0B40),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00920)
);

ninexnine_unit ninexnine_unit_385(
				.clk(clk),
				.rstn(rstn),
				.a0(P0921),
				.a1(P0931),
				.a2(P0941),
				.a3(P0A21),
				.a4(P0A31),
				.a5(P0A41),
				.a6(P0B21),
				.a7(P0B31),
				.a8(P0B41),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01920)
);

ninexnine_unit ninexnine_unit_386(
				.clk(clk),
				.rstn(rstn),
				.a0(P0922),
				.a1(P0932),
				.a2(P0942),
				.a3(P0A22),
				.a4(P0A32),
				.a5(P0A42),
				.a6(P0B22),
				.a7(P0B32),
				.a8(P0B42),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02920)
);

assign C0920=c00920+c01920+c02920;
assign A0920=(C0920>=0)?1:0;

ninexnine_unit ninexnine_unit_387(
				.clk(clk),
				.rstn(rstn),
				.a0(P0930),
				.a1(P0940),
				.a2(P0950),
				.a3(P0A30),
				.a4(P0A40),
				.a5(P0A50),
				.a6(P0B30),
				.a7(P0B40),
				.a8(P0B50),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00930)
);

ninexnine_unit ninexnine_unit_388(
				.clk(clk),
				.rstn(rstn),
				.a0(P0931),
				.a1(P0941),
				.a2(P0951),
				.a3(P0A31),
				.a4(P0A41),
				.a5(P0A51),
				.a6(P0B31),
				.a7(P0B41),
				.a8(P0B51),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01930)
);

ninexnine_unit ninexnine_unit_389(
				.clk(clk),
				.rstn(rstn),
				.a0(P0932),
				.a1(P0942),
				.a2(P0952),
				.a3(P0A32),
				.a4(P0A42),
				.a5(P0A52),
				.a6(P0B32),
				.a7(P0B42),
				.a8(P0B52),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02930)
);

assign C0930=c00930+c01930+c02930;
assign A0930=(C0930>=0)?1:0;

ninexnine_unit ninexnine_unit_390(
				.clk(clk),
				.rstn(rstn),
				.a0(P0940),
				.a1(P0950),
				.a2(P0960),
				.a3(P0A40),
				.a4(P0A50),
				.a5(P0A60),
				.a6(P0B40),
				.a7(P0B50),
				.a8(P0B60),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00940)
);

ninexnine_unit ninexnine_unit_391(
				.clk(clk),
				.rstn(rstn),
				.a0(P0941),
				.a1(P0951),
				.a2(P0961),
				.a3(P0A41),
				.a4(P0A51),
				.a5(P0A61),
				.a6(P0B41),
				.a7(P0B51),
				.a8(P0B61),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01940)
);

ninexnine_unit ninexnine_unit_392(
				.clk(clk),
				.rstn(rstn),
				.a0(P0942),
				.a1(P0952),
				.a2(P0962),
				.a3(P0A42),
				.a4(P0A52),
				.a5(P0A62),
				.a6(P0B42),
				.a7(P0B52),
				.a8(P0B62),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02940)
);

assign C0940=c00940+c01940+c02940;
assign A0940=(C0940>=0)?1:0;

ninexnine_unit ninexnine_unit_393(
				.clk(clk),
				.rstn(rstn),
				.a0(P0950),
				.a1(P0960),
				.a2(P0970),
				.a3(P0A50),
				.a4(P0A60),
				.a5(P0A70),
				.a6(P0B50),
				.a7(P0B60),
				.a8(P0B70),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00950)
);

ninexnine_unit ninexnine_unit_394(
				.clk(clk),
				.rstn(rstn),
				.a0(P0951),
				.a1(P0961),
				.a2(P0971),
				.a3(P0A51),
				.a4(P0A61),
				.a5(P0A71),
				.a6(P0B51),
				.a7(P0B61),
				.a8(P0B71),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01950)
);

ninexnine_unit ninexnine_unit_395(
				.clk(clk),
				.rstn(rstn),
				.a0(P0952),
				.a1(P0962),
				.a2(P0972),
				.a3(P0A52),
				.a4(P0A62),
				.a5(P0A72),
				.a6(P0B52),
				.a7(P0B62),
				.a8(P0B72),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02950)
);

assign C0950=c00950+c01950+c02950;
assign A0950=(C0950>=0)?1:0;

ninexnine_unit ninexnine_unit_396(
				.clk(clk),
				.rstn(rstn),
				.a0(P0960),
				.a1(P0970),
				.a2(P0980),
				.a3(P0A60),
				.a4(P0A70),
				.a5(P0A80),
				.a6(P0B60),
				.a7(P0B70),
				.a8(P0B80),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00960)
);

ninexnine_unit ninexnine_unit_397(
				.clk(clk),
				.rstn(rstn),
				.a0(P0961),
				.a1(P0971),
				.a2(P0981),
				.a3(P0A61),
				.a4(P0A71),
				.a5(P0A81),
				.a6(P0B61),
				.a7(P0B71),
				.a8(P0B81),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01960)
);

ninexnine_unit ninexnine_unit_398(
				.clk(clk),
				.rstn(rstn),
				.a0(P0962),
				.a1(P0972),
				.a2(P0982),
				.a3(P0A62),
				.a4(P0A72),
				.a5(P0A82),
				.a6(P0B62),
				.a7(P0B72),
				.a8(P0B82),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02960)
);

assign C0960=c00960+c01960+c02960;
assign A0960=(C0960>=0)?1:0;

ninexnine_unit ninexnine_unit_399(
				.clk(clk),
				.rstn(rstn),
				.a0(P0970),
				.a1(P0980),
				.a2(P0990),
				.a3(P0A70),
				.a4(P0A80),
				.a5(P0A90),
				.a6(P0B70),
				.a7(P0B80),
				.a8(P0B90),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00970)
);

ninexnine_unit ninexnine_unit_400(
				.clk(clk),
				.rstn(rstn),
				.a0(P0971),
				.a1(P0981),
				.a2(P0991),
				.a3(P0A71),
				.a4(P0A81),
				.a5(P0A91),
				.a6(P0B71),
				.a7(P0B81),
				.a8(P0B91),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01970)
);

ninexnine_unit ninexnine_unit_401(
				.clk(clk),
				.rstn(rstn),
				.a0(P0972),
				.a1(P0982),
				.a2(P0992),
				.a3(P0A72),
				.a4(P0A82),
				.a5(P0A92),
				.a6(P0B72),
				.a7(P0B82),
				.a8(P0B92),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02970)
);

assign C0970=c00970+c01970+c02970;
assign A0970=(C0970>=0)?1:0;

ninexnine_unit ninexnine_unit_402(
				.clk(clk),
				.rstn(rstn),
				.a0(P0980),
				.a1(P0990),
				.a2(P09A0),
				.a3(P0A80),
				.a4(P0A90),
				.a5(P0AA0),
				.a6(P0B80),
				.a7(P0B90),
				.a8(P0BA0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00980)
);

ninexnine_unit ninexnine_unit_403(
				.clk(clk),
				.rstn(rstn),
				.a0(P0981),
				.a1(P0991),
				.a2(P09A1),
				.a3(P0A81),
				.a4(P0A91),
				.a5(P0AA1),
				.a6(P0B81),
				.a7(P0B91),
				.a8(P0BA1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01980)
);

ninexnine_unit ninexnine_unit_404(
				.clk(clk),
				.rstn(rstn),
				.a0(P0982),
				.a1(P0992),
				.a2(P09A2),
				.a3(P0A82),
				.a4(P0A92),
				.a5(P0AA2),
				.a6(P0B82),
				.a7(P0B92),
				.a8(P0BA2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02980)
);

assign C0980=c00980+c01980+c02980;
assign A0980=(C0980>=0)?1:0;

ninexnine_unit ninexnine_unit_405(
				.clk(clk),
				.rstn(rstn),
				.a0(P0990),
				.a1(P09A0),
				.a2(P09B0),
				.a3(P0A90),
				.a4(P0AA0),
				.a5(P0AB0),
				.a6(P0B90),
				.a7(P0BA0),
				.a8(P0BB0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00990)
);

ninexnine_unit ninexnine_unit_406(
				.clk(clk),
				.rstn(rstn),
				.a0(P0991),
				.a1(P09A1),
				.a2(P09B1),
				.a3(P0A91),
				.a4(P0AA1),
				.a5(P0AB1),
				.a6(P0B91),
				.a7(P0BA1),
				.a8(P0BB1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01990)
);

ninexnine_unit ninexnine_unit_407(
				.clk(clk),
				.rstn(rstn),
				.a0(P0992),
				.a1(P09A2),
				.a2(P09B2),
				.a3(P0A92),
				.a4(P0AA2),
				.a5(P0AB2),
				.a6(P0B92),
				.a7(P0BA2),
				.a8(P0BB2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02990)
);

assign C0990=c00990+c01990+c02990;
assign A0990=(C0990>=0)?1:0;

ninexnine_unit ninexnine_unit_408(
				.clk(clk),
				.rstn(rstn),
				.a0(P09A0),
				.a1(P09B0),
				.a2(P09C0),
				.a3(P0AA0),
				.a4(P0AB0),
				.a5(P0AC0),
				.a6(P0BA0),
				.a7(P0BB0),
				.a8(P0BC0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c009A0)
);

ninexnine_unit ninexnine_unit_409(
				.clk(clk),
				.rstn(rstn),
				.a0(P09A1),
				.a1(P09B1),
				.a2(P09C1),
				.a3(P0AA1),
				.a4(P0AB1),
				.a5(P0AC1),
				.a6(P0BA1),
				.a7(P0BB1),
				.a8(P0BC1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c019A0)
);

ninexnine_unit ninexnine_unit_410(
				.clk(clk),
				.rstn(rstn),
				.a0(P09A2),
				.a1(P09B2),
				.a2(P09C2),
				.a3(P0AA2),
				.a4(P0AB2),
				.a5(P0AC2),
				.a6(P0BA2),
				.a7(P0BB2),
				.a8(P0BC2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c029A0)
);

assign C09A0=c009A0+c019A0+c029A0;
assign A09A0=(C09A0>=0)?1:0;

ninexnine_unit ninexnine_unit_411(
				.clk(clk),
				.rstn(rstn),
				.a0(P09B0),
				.a1(P09C0),
				.a2(P09D0),
				.a3(P0AB0),
				.a4(P0AC0),
				.a5(P0AD0),
				.a6(P0BB0),
				.a7(P0BC0),
				.a8(P0BD0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c009B0)
);

ninexnine_unit ninexnine_unit_412(
				.clk(clk),
				.rstn(rstn),
				.a0(P09B1),
				.a1(P09C1),
				.a2(P09D1),
				.a3(P0AB1),
				.a4(P0AC1),
				.a5(P0AD1),
				.a6(P0BB1),
				.a7(P0BC1),
				.a8(P0BD1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c019B0)
);

ninexnine_unit ninexnine_unit_413(
				.clk(clk),
				.rstn(rstn),
				.a0(P09B2),
				.a1(P09C2),
				.a2(P09D2),
				.a3(P0AB2),
				.a4(P0AC2),
				.a5(P0AD2),
				.a6(P0BB2),
				.a7(P0BC2),
				.a8(P0BD2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c029B0)
);

assign C09B0=c009B0+c019B0+c029B0;
assign A09B0=(C09B0>=0)?1:0;

ninexnine_unit ninexnine_unit_414(
				.clk(clk),
				.rstn(rstn),
				.a0(P09C0),
				.a1(P09D0),
				.a2(P09E0),
				.a3(P0AC0),
				.a4(P0AD0),
				.a5(P0AE0),
				.a6(P0BC0),
				.a7(P0BD0),
				.a8(P0BE0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c009C0)
);

ninexnine_unit ninexnine_unit_415(
				.clk(clk),
				.rstn(rstn),
				.a0(P09C1),
				.a1(P09D1),
				.a2(P09E1),
				.a3(P0AC1),
				.a4(P0AD1),
				.a5(P0AE1),
				.a6(P0BC1),
				.a7(P0BD1),
				.a8(P0BE1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c019C0)
);

ninexnine_unit ninexnine_unit_416(
				.clk(clk),
				.rstn(rstn),
				.a0(P09C2),
				.a1(P09D2),
				.a2(P09E2),
				.a3(P0AC2),
				.a4(P0AD2),
				.a5(P0AE2),
				.a6(P0BC2),
				.a7(P0BD2),
				.a8(P0BE2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c029C0)
);

assign C09C0=c009C0+c019C0+c029C0;
assign A09C0=(C09C0>=0)?1:0;

ninexnine_unit ninexnine_unit_417(
				.clk(clk),
				.rstn(rstn),
				.a0(P09D0),
				.a1(P09E0),
				.a2(P09F0),
				.a3(P0AD0),
				.a4(P0AE0),
				.a5(P0AF0),
				.a6(P0BD0),
				.a7(P0BE0),
				.a8(P0BF0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c009D0)
);

ninexnine_unit ninexnine_unit_418(
				.clk(clk),
				.rstn(rstn),
				.a0(P09D1),
				.a1(P09E1),
				.a2(P09F1),
				.a3(P0AD1),
				.a4(P0AE1),
				.a5(P0AF1),
				.a6(P0BD1),
				.a7(P0BE1),
				.a8(P0BF1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c019D0)
);

ninexnine_unit ninexnine_unit_419(
				.clk(clk),
				.rstn(rstn),
				.a0(P09D2),
				.a1(P09E2),
				.a2(P09F2),
				.a3(P0AD2),
				.a4(P0AE2),
				.a5(P0AF2),
				.a6(P0BD2),
				.a7(P0BE2),
				.a8(P0BF2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c029D0)
);

assign C09D0=c009D0+c019D0+c029D0;
assign A09D0=(C09D0>=0)?1:0;

ninexnine_unit ninexnine_unit_420(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A00),
				.a1(P0A10),
				.a2(P0A20),
				.a3(P0B00),
				.a4(P0B10),
				.a5(P0B20),
				.a6(P0C00),
				.a7(P0C10),
				.a8(P0C20),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00A00)
);

ninexnine_unit ninexnine_unit_421(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A01),
				.a1(P0A11),
				.a2(P0A21),
				.a3(P0B01),
				.a4(P0B11),
				.a5(P0B21),
				.a6(P0C01),
				.a7(P0C11),
				.a8(P0C21),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01A00)
);

ninexnine_unit ninexnine_unit_422(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A02),
				.a1(P0A12),
				.a2(P0A22),
				.a3(P0B02),
				.a4(P0B12),
				.a5(P0B22),
				.a6(P0C02),
				.a7(P0C12),
				.a8(P0C22),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02A00)
);

assign C0A00=c00A00+c01A00+c02A00;
assign A0A00=(C0A00>=0)?1:0;

ninexnine_unit ninexnine_unit_423(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A10),
				.a1(P0A20),
				.a2(P0A30),
				.a3(P0B10),
				.a4(P0B20),
				.a5(P0B30),
				.a6(P0C10),
				.a7(P0C20),
				.a8(P0C30),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00A10)
);

ninexnine_unit ninexnine_unit_424(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A11),
				.a1(P0A21),
				.a2(P0A31),
				.a3(P0B11),
				.a4(P0B21),
				.a5(P0B31),
				.a6(P0C11),
				.a7(P0C21),
				.a8(P0C31),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01A10)
);

ninexnine_unit ninexnine_unit_425(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A12),
				.a1(P0A22),
				.a2(P0A32),
				.a3(P0B12),
				.a4(P0B22),
				.a5(P0B32),
				.a6(P0C12),
				.a7(P0C22),
				.a8(P0C32),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02A10)
);

assign C0A10=c00A10+c01A10+c02A10;
assign A0A10=(C0A10>=0)?1:0;

ninexnine_unit ninexnine_unit_426(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A20),
				.a1(P0A30),
				.a2(P0A40),
				.a3(P0B20),
				.a4(P0B30),
				.a5(P0B40),
				.a6(P0C20),
				.a7(P0C30),
				.a8(P0C40),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00A20)
);

ninexnine_unit ninexnine_unit_427(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A21),
				.a1(P0A31),
				.a2(P0A41),
				.a3(P0B21),
				.a4(P0B31),
				.a5(P0B41),
				.a6(P0C21),
				.a7(P0C31),
				.a8(P0C41),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01A20)
);

ninexnine_unit ninexnine_unit_428(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A22),
				.a1(P0A32),
				.a2(P0A42),
				.a3(P0B22),
				.a4(P0B32),
				.a5(P0B42),
				.a6(P0C22),
				.a7(P0C32),
				.a8(P0C42),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02A20)
);

assign C0A20=c00A20+c01A20+c02A20;
assign A0A20=(C0A20>=0)?1:0;

ninexnine_unit ninexnine_unit_429(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A30),
				.a1(P0A40),
				.a2(P0A50),
				.a3(P0B30),
				.a4(P0B40),
				.a5(P0B50),
				.a6(P0C30),
				.a7(P0C40),
				.a8(P0C50),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00A30)
);

ninexnine_unit ninexnine_unit_430(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A31),
				.a1(P0A41),
				.a2(P0A51),
				.a3(P0B31),
				.a4(P0B41),
				.a5(P0B51),
				.a6(P0C31),
				.a7(P0C41),
				.a8(P0C51),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01A30)
);

ninexnine_unit ninexnine_unit_431(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A32),
				.a1(P0A42),
				.a2(P0A52),
				.a3(P0B32),
				.a4(P0B42),
				.a5(P0B52),
				.a6(P0C32),
				.a7(P0C42),
				.a8(P0C52),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02A30)
);

assign C0A30=c00A30+c01A30+c02A30;
assign A0A30=(C0A30>=0)?1:0;

ninexnine_unit ninexnine_unit_432(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A40),
				.a1(P0A50),
				.a2(P0A60),
				.a3(P0B40),
				.a4(P0B50),
				.a5(P0B60),
				.a6(P0C40),
				.a7(P0C50),
				.a8(P0C60),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00A40)
);

ninexnine_unit ninexnine_unit_433(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A41),
				.a1(P0A51),
				.a2(P0A61),
				.a3(P0B41),
				.a4(P0B51),
				.a5(P0B61),
				.a6(P0C41),
				.a7(P0C51),
				.a8(P0C61),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01A40)
);

ninexnine_unit ninexnine_unit_434(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A42),
				.a1(P0A52),
				.a2(P0A62),
				.a3(P0B42),
				.a4(P0B52),
				.a5(P0B62),
				.a6(P0C42),
				.a7(P0C52),
				.a8(P0C62),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02A40)
);

assign C0A40=c00A40+c01A40+c02A40;
assign A0A40=(C0A40>=0)?1:0;

ninexnine_unit ninexnine_unit_435(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A50),
				.a1(P0A60),
				.a2(P0A70),
				.a3(P0B50),
				.a4(P0B60),
				.a5(P0B70),
				.a6(P0C50),
				.a7(P0C60),
				.a8(P0C70),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00A50)
);

ninexnine_unit ninexnine_unit_436(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A51),
				.a1(P0A61),
				.a2(P0A71),
				.a3(P0B51),
				.a4(P0B61),
				.a5(P0B71),
				.a6(P0C51),
				.a7(P0C61),
				.a8(P0C71),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01A50)
);

ninexnine_unit ninexnine_unit_437(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A52),
				.a1(P0A62),
				.a2(P0A72),
				.a3(P0B52),
				.a4(P0B62),
				.a5(P0B72),
				.a6(P0C52),
				.a7(P0C62),
				.a8(P0C72),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02A50)
);

assign C0A50=c00A50+c01A50+c02A50;
assign A0A50=(C0A50>=0)?1:0;

ninexnine_unit ninexnine_unit_438(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A60),
				.a1(P0A70),
				.a2(P0A80),
				.a3(P0B60),
				.a4(P0B70),
				.a5(P0B80),
				.a6(P0C60),
				.a7(P0C70),
				.a8(P0C80),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00A60)
);

ninexnine_unit ninexnine_unit_439(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A61),
				.a1(P0A71),
				.a2(P0A81),
				.a3(P0B61),
				.a4(P0B71),
				.a5(P0B81),
				.a6(P0C61),
				.a7(P0C71),
				.a8(P0C81),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01A60)
);

ninexnine_unit ninexnine_unit_440(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A62),
				.a1(P0A72),
				.a2(P0A82),
				.a3(P0B62),
				.a4(P0B72),
				.a5(P0B82),
				.a6(P0C62),
				.a7(P0C72),
				.a8(P0C82),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02A60)
);

assign C0A60=c00A60+c01A60+c02A60;
assign A0A60=(C0A60>=0)?1:0;

ninexnine_unit ninexnine_unit_441(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A70),
				.a1(P0A80),
				.a2(P0A90),
				.a3(P0B70),
				.a4(P0B80),
				.a5(P0B90),
				.a6(P0C70),
				.a7(P0C80),
				.a8(P0C90),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00A70)
);

ninexnine_unit ninexnine_unit_442(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A71),
				.a1(P0A81),
				.a2(P0A91),
				.a3(P0B71),
				.a4(P0B81),
				.a5(P0B91),
				.a6(P0C71),
				.a7(P0C81),
				.a8(P0C91),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01A70)
);

ninexnine_unit ninexnine_unit_443(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A72),
				.a1(P0A82),
				.a2(P0A92),
				.a3(P0B72),
				.a4(P0B82),
				.a5(P0B92),
				.a6(P0C72),
				.a7(P0C82),
				.a8(P0C92),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02A70)
);

assign C0A70=c00A70+c01A70+c02A70;
assign A0A70=(C0A70>=0)?1:0;

ninexnine_unit ninexnine_unit_444(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A80),
				.a1(P0A90),
				.a2(P0AA0),
				.a3(P0B80),
				.a4(P0B90),
				.a5(P0BA0),
				.a6(P0C80),
				.a7(P0C90),
				.a8(P0CA0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00A80)
);

ninexnine_unit ninexnine_unit_445(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A81),
				.a1(P0A91),
				.a2(P0AA1),
				.a3(P0B81),
				.a4(P0B91),
				.a5(P0BA1),
				.a6(P0C81),
				.a7(P0C91),
				.a8(P0CA1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01A80)
);

ninexnine_unit ninexnine_unit_446(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A82),
				.a1(P0A92),
				.a2(P0AA2),
				.a3(P0B82),
				.a4(P0B92),
				.a5(P0BA2),
				.a6(P0C82),
				.a7(P0C92),
				.a8(P0CA2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02A80)
);

assign C0A80=c00A80+c01A80+c02A80;
assign A0A80=(C0A80>=0)?1:0;

ninexnine_unit ninexnine_unit_447(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A90),
				.a1(P0AA0),
				.a2(P0AB0),
				.a3(P0B90),
				.a4(P0BA0),
				.a5(P0BB0),
				.a6(P0C90),
				.a7(P0CA0),
				.a8(P0CB0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00A90)
);

ninexnine_unit ninexnine_unit_448(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A91),
				.a1(P0AA1),
				.a2(P0AB1),
				.a3(P0B91),
				.a4(P0BA1),
				.a5(P0BB1),
				.a6(P0C91),
				.a7(P0CA1),
				.a8(P0CB1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01A90)
);

ninexnine_unit ninexnine_unit_449(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A92),
				.a1(P0AA2),
				.a2(P0AB2),
				.a3(P0B92),
				.a4(P0BA2),
				.a5(P0BB2),
				.a6(P0C92),
				.a7(P0CA2),
				.a8(P0CB2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02A90)
);

assign C0A90=c00A90+c01A90+c02A90;
assign A0A90=(C0A90>=0)?1:0;

ninexnine_unit ninexnine_unit_450(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AA0),
				.a1(P0AB0),
				.a2(P0AC0),
				.a3(P0BA0),
				.a4(P0BB0),
				.a5(P0BC0),
				.a6(P0CA0),
				.a7(P0CB0),
				.a8(P0CC0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00AA0)
);

ninexnine_unit ninexnine_unit_451(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AA1),
				.a1(P0AB1),
				.a2(P0AC1),
				.a3(P0BA1),
				.a4(P0BB1),
				.a5(P0BC1),
				.a6(P0CA1),
				.a7(P0CB1),
				.a8(P0CC1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01AA0)
);

ninexnine_unit ninexnine_unit_452(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AA2),
				.a1(P0AB2),
				.a2(P0AC2),
				.a3(P0BA2),
				.a4(P0BB2),
				.a5(P0BC2),
				.a6(P0CA2),
				.a7(P0CB2),
				.a8(P0CC2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02AA0)
);

assign C0AA0=c00AA0+c01AA0+c02AA0;
assign A0AA0=(C0AA0>=0)?1:0;

ninexnine_unit ninexnine_unit_453(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AB0),
				.a1(P0AC0),
				.a2(P0AD0),
				.a3(P0BB0),
				.a4(P0BC0),
				.a5(P0BD0),
				.a6(P0CB0),
				.a7(P0CC0),
				.a8(P0CD0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00AB0)
);

ninexnine_unit ninexnine_unit_454(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AB1),
				.a1(P0AC1),
				.a2(P0AD1),
				.a3(P0BB1),
				.a4(P0BC1),
				.a5(P0BD1),
				.a6(P0CB1),
				.a7(P0CC1),
				.a8(P0CD1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01AB0)
);

ninexnine_unit ninexnine_unit_455(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AB2),
				.a1(P0AC2),
				.a2(P0AD2),
				.a3(P0BB2),
				.a4(P0BC2),
				.a5(P0BD2),
				.a6(P0CB2),
				.a7(P0CC2),
				.a8(P0CD2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02AB0)
);

assign C0AB0=c00AB0+c01AB0+c02AB0;
assign A0AB0=(C0AB0>=0)?1:0;

ninexnine_unit ninexnine_unit_456(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AC0),
				.a1(P0AD0),
				.a2(P0AE0),
				.a3(P0BC0),
				.a4(P0BD0),
				.a5(P0BE0),
				.a6(P0CC0),
				.a7(P0CD0),
				.a8(P0CE0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00AC0)
);

ninexnine_unit ninexnine_unit_457(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AC1),
				.a1(P0AD1),
				.a2(P0AE1),
				.a3(P0BC1),
				.a4(P0BD1),
				.a5(P0BE1),
				.a6(P0CC1),
				.a7(P0CD1),
				.a8(P0CE1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01AC0)
);

ninexnine_unit ninexnine_unit_458(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AC2),
				.a1(P0AD2),
				.a2(P0AE2),
				.a3(P0BC2),
				.a4(P0BD2),
				.a5(P0BE2),
				.a6(P0CC2),
				.a7(P0CD2),
				.a8(P0CE2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02AC0)
);

assign C0AC0=c00AC0+c01AC0+c02AC0;
assign A0AC0=(C0AC0>=0)?1:0;

ninexnine_unit ninexnine_unit_459(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AD0),
				.a1(P0AE0),
				.a2(P0AF0),
				.a3(P0BD0),
				.a4(P0BE0),
				.a5(P0BF0),
				.a6(P0CD0),
				.a7(P0CE0),
				.a8(P0CF0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00AD0)
);

ninexnine_unit ninexnine_unit_460(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AD1),
				.a1(P0AE1),
				.a2(P0AF1),
				.a3(P0BD1),
				.a4(P0BE1),
				.a5(P0BF1),
				.a6(P0CD1),
				.a7(P0CE1),
				.a8(P0CF1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01AD0)
);

ninexnine_unit ninexnine_unit_461(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AD2),
				.a1(P0AE2),
				.a2(P0AF2),
				.a3(P0BD2),
				.a4(P0BE2),
				.a5(P0BF2),
				.a6(P0CD2),
				.a7(P0CE2),
				.a8(P0CF2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02AD0)
);

assign C0AD0=c00AD0+c01AD0+c02AD0;
assign A0AD0=(C0AD0>=0)?1:0;

ninexnine_unit ninexnine_unit_462(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B00),
				.a1(P0B10),
				.a2(P0B20),
				.a3(P0C00),
				.a4(P0C10),
				.a5(P0C20),
				.a6(P0D00),
				.a7(P0D10),
				.a8(P0D20),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00B00)
);

ninexnine_unit ninexnine_unit_463(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B01),
				.a1(P0B11),
				.a2(P0B21),
				.a3(P0C01),
				.a4(P0C11),
				.a5(P0C21),
				.a6(P0D01),
				.a7(P0D11),
				.a8(P0D21),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01B00)
);

ninexnine_unit ninexnine_unit_464(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B02),
				.a1(P0B12),
				.a2(P0B22),
				.a3(P0C02),
				.a4(P0C12),
				.a5(P0C22),
				.a6(P0D02),
				.a7(P0D12),
				.a8(P0D22),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02B00)
);

assign C0B00=c00B00+c01B00+c02B00;
assign A0B00=(C0B00>=0)?1:0;

ninexnine_unit ninexnine_unit_465(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B10),
				.a1(P0B20),
				.a2(P0B30),
				.a3(P0C10),
				.a4(P0C20),
				.a5(P0C30),
				.a6(P0D10),
				.a7(P0D20),
				.a8(P0D30),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00B10)
);

ninexnine_unit ninexnine_unit_466(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B11),
				.a1(P0B21),
				.a2(P0B31),
				.a3(P0C11),
				.a4(P0C21),
				.a5(P0C31),
				.a6(P0D11),
				.a7(P0D21),
				.a8(P0D31),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01B10)
);

ninexnine_unit ninexnine_unit_467(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B12),
				.a1(P0B22),
				.a2(P0B32),
				.a3(P0C12),
				.a4(P0C22),
				.a5(P0C32),
				.a6(P0D12),
				.a7(P0D22),
				.a8(P0D32),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02B10)
);

assign C0B10=c00B10+c01B10+c02B10;
assign A0B10=(C0B10>=0)?1:0;

ninexnine_unit ninexnine_unit_468(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B20),
				.a1(P0B30),
				.a2(P0B40),
				.a3(P0C20),
				.a4(P0C30),
				.a5(P0C40),
				.a6(P0D20),
				.a7(P0D30),
				.a8(P0D40),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00B20)
);

ninexnine_unit ninexnine_unit_469(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B21),
				.a1(P0B31),
				.a2(P0B41),
				.a3(P0C21),
				.a4(P0C31),
				.a5(P0C41),
				.a6(P0D21),
				.a7(P0D31),
				.a8(P0D41),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01B20)
);

ninexnine_unit ninexnine_unit_470(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B22),
				.a1(P0B32),
				.a2(P0B42),
				.a3(P0C22),
				.a4(P0C32),
				.a5(P0C42),
				.a6(P0D22),
				.a7(P0D32),
				.a8(P0D42),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02B20)
);

assign C0B20=c00B20+c01B20+c02B20;
assign A0B20=(C0B20>=0)?1:0;

ninexnine_unit ninexnine_unit_471(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B30),
				.a1(P0B40),
				.a2(P0B50),
				.a3(P0C30),
				.a4(P0C40),
				.a5(P0C50),
				.a6(P0D30),
				.a7(P0D40),
				.a8(P0D50),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00B30)
);

ninexnine_unit ninexnine_unit_472(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B31),
				.a1(P0B41),
				.a2(P0B51),
				.a3(P0C31),
				.a4(P0C41),
				.a5(P0C51),
				.a6(P0D31),
				.a7(P0D41),
				.a8(P0D51),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01B30)
);

ninexnine_unit ninexnine_unit_473(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B32),
				.a1(P0B42),
				.a2(P0B52),
				.a3(P0C32),
				.a4(P0C42),
				.a5(P0C52),
				.a6(P0D32),
				.a7(P0D42),
				.a8(P0D52),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02B30)
);

assign C0B30=c00B30+c01B30+c02B30;
assign A0B30=(C0B30>=0)?1:0;

ninexnine_unit ninexnine_unit_474(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B40),
				.a1(P0B50),
				.a2(P0B60),
				.a3(P0C40),
				.a4(P0C50),
				.a5(P0C60),
				.a6(P0D40),
				.a7(P0D50),
				.a8(P0D60),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00B40)
);

ninexnine_unit ninexnine_unit_475(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B41),
				.a1(P0B51),
				.a2(P0B61),
				.a3(P0C41),
				.a4(P0C51),
				.a5(P0C61),
				.a6(P0D41),
				.a7(P0D51),
				.a8(P0D61),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01B40)
);

ninexnine_unit ninexnine_unit_476(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B42),
				.a1(P0B52),
				.a2(P0B62),
				.a3(P0C42),
				.a4(P0C52),
				.a5(P0C62),
				.a6(P0D42),
				.a7(P0D52),
				.a8(P0D62),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02B40)
);

assign C0B40=c00B40+c01B40+c02B40;
assign A0B40=(C0B40>=0)?1:0;

ninexnine_unit ninexnine_unit_477(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B50),
				.a1(P0B60),
				.a2(P0B70),
				.a3(P0C50),
				.a4(P0C60),
				.a5(P0C70),
				.a6(P0D50),
				.a7(P0D60),
				.a8(P0D70),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00B50)
);

ninexnine_unit ninexnine_unit_478(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B51),
				.a1(P0B61),
				.a2(P0B71),
				.a3(P0C51),
				.a4(P0C61),
				.a5(P0C71),
				.a6(P0D51),
				.a7(P0D61),
				.a8(P0D71),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01B50)
);

ninexnine_unit ninexnine_unit_479(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B52),
				.a1(P0B62),
				.a2(P0B72),
				.a3(P0C52),
				.a4(P0C62),
				.a5(P0C72),
				.a6(P0D52),
				.a7(P0D62),
				.a8(P0D72),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02B50)
);

assign C0B50=c00B50+c01B50+c02B50;
assign A0B50=(C0B50>=0)?1:0;

ninexnine_unit ninexnine_unit_480(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B60),
				.a1(P0B70),
				.a2(P0B80),
				.a3(P0C60),
				.a4(P0C70),
				.a5(P0C80),
				.a6(P0D60),
				.a7(P0D70),
				.a8(P0D80),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00B60)
);

ninexnine_unit ninexnine_unit_481(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B61),
				.a1(P0B71),
				.a2(P0B81),
				.a3(P0C61),
				.a4(P0C71),
				.a5(P0C81),
				.a6(P0D61),
				.a7(P0D71),
				.a8(P0D81),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01B60)
);

ninexnine_unit ninexnine_unit_482(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B62),
				.a1(P0B72),
				.a2(P0B82),
				.a3(P0C62),
				.a4(P0C72),
				.a5(P0C82),
				.a6(P0D62),
				.a7(P0D72),
				.a8(P0D82),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02B60)
);

assign C0B60=c00B60+c01B60+c02B60;
assign A0B60=(C0B60>=0)?1:0;

ninexnine_unit ninexnine_unit_483(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B70),
				.a1(P0B80),
				.a2(P0B90),
				.a3(P0C70),
				.a4(P0C80),
				.a5(P0C90),
				.a6(P0D70),
				.a7(P0D80),
				.a8(P0D90),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00B70)
);

ninexnine_unit ninexnine_unit_484(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B71),
				.a1(P0B81),
				.a2(P0B91),
				.a3(P0C71),
				.a4(P0C81),
				.a5(P0C91),
				.a6(P0D71),
				.a7(P0D81),
				.a8(P0D91),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01B70)
);

ninexnine_unit ninexnine_unit_485(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B72),
				.a1(P0B82),
				.a2(P0B92),
				.a3(P0C72),
				.a4(P0C82),
				.a5(P0C92),
				.a6(P0D72),
				.a7(P0D82),
				.a8(P0D92),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02B70)
);

assign C0B70=c00B70+c01B70+c02B70;
assign A0B70=(C0B70>=0)?1:0;

ninexnine_unit ninexnine_unit_486(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B80),
				.a1(P0B90),
				.a2(P0BA0),
				.a3(P0C80),
				.a4(P0C90),
				.a5(P0CA0),
				.a6(P0D80),
				.a7(P0D90),
				.a8(P0DA0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00B80)
);

ninexnine_unit ninexnine_unit_487(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B81),
				.a1(P0B91),
				.a2(P0BA1),
				.a3(P0C81),
				.a4(P0C91),
				.a5(P0CA1),
				.a6(P0D81),
				.a7(P0D91),
				.a8(P0DA1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01B80)
);

ninexnine_unit ninexnine_unit_488(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B82),
				.a1(P0B92),
				.a2(P0BA2),
				.a3(P0C82),
				.a4(P0C92),
				.a5(P0CA2),
				.a6(P0D82),
				.a7(P0D92),
				.a8(P0DA2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02B80)
);

assign C0B80=c00B80+c01B80+c02B80;
assign A0B80=(C0B80>=0)?1:0;

ninexnine_unit ninexnine_unit_489(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B90),
				.a1(P0BA0),
				.a2(P0BB0),
				.a3(P0C90),
				.a4(P0CA0),
				.a5(P0CB0),
				.a6(P0D90),
				.a7(P0DA0),
				.a8(P0DB0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00B90)
);

ninexnine_unit ninexnine_unit_490(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B91),
				.a1(P0BA1),
				.a2(P0BB1),
				.a3(P0C91),
				.a4(P0CA1),
				.a5(P0CB1),
				.a6(P0D91),
				.a7(P0DA1),
				.a8(P0DB1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01B90)
);

ninexnine_unit ninexnine_unit_491(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B92),
				.a1(P0BA2),
				.a2(P0BB2),
				.a3(P0C92),
				.a4(P0CA2),
				.a5(P0CB2),
				.a6(P0D92),
				.a7(P0DA2),
				.a8(P0DB2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02B90)
);

assign C0B90=c00B90+c01B90+c02B90;
assign A0B90=(C0B90>=0)?1:0;

ninexnine_unit ninexnine_unit_492(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BA0),
				.a1(P0BB0),
				.a2(P0BC0),
				.a3(P0CA0),
				.a4(P0CB0),
				.a5(P0CC0),
				.a6(P0DA0),
				.a7(P0DB0),
				.a8(P0DC0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00BA0)
);

ninexnine_unit ninexnine_unit_493(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BA1),
				.a1(P0BB1),
				.a2(P0BC1),
				.a3(P0CA1),
				.a4(P0CB1),
				.a5(P0CC1),
				.a6(P0DA1),
				.a7(P0DB1),
				.a8(P0DC1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01BA0)
);

ninexnine_unit ninexnine_unit_494(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BA2),
				.a1(P0BB2),
				.a2(P0BC2),
				.a3(P0CA2),
				.a4(P0CB2),
				.a5(P0CC2),
				.a6(P0DA2),
				.a7(P0DB2),
				.a8(P0DC2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02BA0)
);

assign C0BA0=c00BA0+c01BA0+c02BA0;
assign A0BA0=(C0BA0>=0)?1:0;

ninexnine_unit ninexnine_unit_495(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BB0),
				.a1(P0BC0),
				.a2(P0BD0),
				.a3(P0CB0),
				.a4(P0CC0),
				.a5(P0CD0),
				.a6(P0DB0),
				.a7(P0DC0),
				.a8(P0DD0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00BB0)
);

ninexnine_unit ninexnine_unit_496(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BB1),
				.a1(P0BC1),
				.a2(P0BD1),
				.a3(P0CB1),
				.a4(P0CC1),
				.a5(P0CD1),
				.a6(P0DB1),
				.a7(P0DC1),
				.a8(P0DD1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01BB0)
);

ninexnine_unit ninexnine_unit_497(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BB2),
				.a1(P0BC2),
				.a2(P0BD2),
				.a3(P0CB2),
				.a4(P0CC2),
				.a5(P0CD2),
				.a6(P0DB2),
				.a7(P0DC2),
				.a8(P0DD2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02BB0)
);

assign C0BB0=c00BB0+c01BB0+c02BB0;
assign A0BB0=(C0BB0>=0)?1:0;

ninexnine_unit ninexnine_unit_498(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BC0),
				.a1(P0BD0),
				.a2(P0BE0),
				.a3(P0CC0),
				.a4(P0CD0),
				.a5(P0CE0),
				.a6(P0DC0),
				.a7(P0DD0),
				.a8(P0DE0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00BC0)
);

ninexnine_unit ninexnine_unit_499(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BC1),
				.a1(P0BD1),
				.a2(P0BE1),
				.a3(P0CC1),
				.a4(P0CD1),
				.a5(P0CE1),
				.a6(P0DC1),
				.a7(P0DD1),
				.a8(P0DE1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01BC0)
);

ninexnine_unit ninexnine_unit_500(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BC2),
				.a1(P0BD2),
				.a2(P0BE2),
				.a3(P0CC2),
				.a4(P0CD2),
				.a5(P0CE2),
				.a6(P0DC2),
				.a7(P0DD2),
				.a8(P0DE2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02BC0)
);

assign C0BC0=c00BC0+c01BC0+c02BC0;
assign A0BC0=(C0BC0>=0)?1:0;

ninexnine_unit ninexnine_unit_501(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BD0),
				.a1(P0BE0),
				.a2(P0BF0),
				.a3(P0CD0),
				.a4(P0CE0),
				.a5(P0CF0),
				.a6(P0DD0),
				.a7(P0DE0),
				.a8(P0DF0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00BD0)
);

ninexnine_unit ninexnine_unit_502(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BD1),
				.a1(P0BE1),
				.a2(P0BF1),
				.a3(P0CD1),
				.a4(P0CE1),
				.a5(P0CF1),
				.a6(P0DD1),
				.a7(P0DE1),
				.a8(P0DF1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01BD0)
);

ninexnine_unit ninexnine_unit_503(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BD2),
				.a1(P0BE2),
				.a2(P0BF2),
				.a3(P0CD2),
				.a4(P0CE2),
				.a5(P0CF2),
				.a6(P0DD2),
				.a7(P0DE2),
				.a8(P0DF2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02BD0)
);

assign C0BD0=c00BD0+c01BD0+c02BD0;
assign A0BD0=(C0BD0>=0)?1:0;

ninexnine_unit ninexnine_unit_504(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C00),
				.a1(P0C10),
				.a2(P0C20),
				.a3(P0D00),
				.a4(P0D10),
				.a5(P0D20),
				.a6(P0E00),
				.a7(P0E10),
				.a8(P0E20),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00C00)
);

ninexnine_unit ninexnine_unit_505(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C01),
				.a1(P0C11),
				.a2(P0C21),
				.a3(P0D01),
				.a4(P0D11),
				.a5(P0D21),
				.a6(P0E01),
				.a7(P0E11),
				.a8(P0E21),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01C00)
);

ninexnine_unit ninexnine_unit_506(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C02),
				.a1(P0C12),
				.a2(P0C22),
				.a3(P0D02),
				.a4(P0D12),
				.a5(P0D22),
				.a6(P0E02),
				.a7(P0E12),
				.a8(P0E22),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02C00)
);

assign C0C00=c00C00+c01C00+c02C00;
assign A0C00=(C0C00>=0)?1:0;

ninexnine_unit ninexnine_unit_507(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C10),
				.a1(P0C20),
				.a2(P0C30),
				.a3(P0D10),
				.a4(P0D20),
				.a5(P0D30),
				.a6(P0E10),
				.a7(P0E20),
				.a8(P0E30),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00C10)
);

ninexnine_unit ninexnine_unit_508(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C11),
				.a1(P0C21),
				.a2(P0C31),
				.a3(P0D11),
				.a4(P0D21),
				.a5(P0D31),
				.a6(P0E11),
				.a7(P0E21),
				.a8(P0E31),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01C10)
);

ninexnine_unit ninexnine_unit_509(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C12),
				.a1(P0C22),
				.a2(P0C32),
				.a3(P0D12),
				.a4(P0D22),
				.a5(P0D32),
				.a6(P0E12),
				.a7(P0E22),
				.a8(P0E32),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02C10)
);

assign C0C10=c00C10+c01C10+c02C10;
assign A0C10=(C0C10>=0)?1:0;

ninexnine_unit ninexnine_unit_510(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C20),
				.a1(P0C30),
				.a2(P0C40),
				.a3(P0D20),
				.a4(P0D30),
				.a5(P0D40),
				.a6(P0E20),
				.a7(P0E30),
				.a8(P0E40),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00C20)
);

ninexnine_unit ninexnine_unit_511(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C21),
				.a1(P0C31),
				.a2(P0C41),
				.a3(P0D21),
				.a4(P0D31),
				.a5(P0D41),
				.a6(P0E21),
				.a7(P0E31),
				.a8(P0E41),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01C20)
);

ninexnine_unit ninexnine_unit_512(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C22),
				.a1(P0C32),
				.a2(P0C42),
				.a3(P0D22),
				.a4(P0D32),
				.a5(P0D42),
				.a6(P0E22),
				.a7(P0E32),
				.a8(P0E42),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02C20)
);

assign C0C20=c00C20+c01C20+c02C20;
assign A0C20=(C0C20>=0)?1:0;

ninexnine_unit ninexnine_unit_513(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C30),
				.a1(P0C40),
				.a2(P0C50),
				.a3(P0D30),
				.a4(P0D40),
				.a5(P0D50),
				.a6(P0E30),
				.a7(P0E40),
				.a8(P0E50),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00C30)
);

ninexnine_unit ninexnine_unit_514(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C31),
				.a1(P0C41),
				.a2(P0C51),
				.a3(P0D31),
				.a4(P0D41),
				.a5(P0D51),
				.a6(P0E31),
				.a7(P0E41),
				.a8(P0E51),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01C30)
);

ninexnine_unit ninexnine_unit_515(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C32),
				.a1(P0C42),
				.a2(P0C52),
				.a3(P0D32),
				.a4(P0D42),
				.a5(P0D52),
				.a6(P0E32),
				.a7(P0E42),
				.a8(P0E52),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02C30)
);

assign C0C30=c00C30+c01C30+c02C30;
assign A0C30=(C0C30>=0)?1:0;

ninexnine_unit ninexnine_unit_516(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C40),
				.a1(P0C50),
				.a2(P0C60),
				.a3(P0D40),
				.a4(P0D50),
				.a5(P0D60),
				.a6(P0E40),
				.a7(P0E50),
				.a8(P0E60),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00C40)
);

ninexnine_unit ninexnine_unit_517(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C41),
				.a1(P0C51),
				.a2(P0C61),
				.a3(P0D41),
				.a4(P0D51),
				.a5(P0D61),
				.a6(P0E41),
				.a7(P0E51),
				.a8(P0E61),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01C40)
);

ninexnine_unit ninexnine_unit_518(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C42),
				.a1(P0C52),
				.a2(P0C62),
				.a3(P0D42),
				.a4(P0D52),
				.a5(P0D62),
				.a6(P0E42),
				.a7(P0E52),
				.a8(P0E62),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02C40)
);

assign C0C40=c00C40+c01C40+c02C40;
assign A0C40=(C0C40>=0)?1:0;

ninexnine_unit ninexnine_unit_519(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C50),
				.a1(P0C60),
				.a2(P0C70),
				.a3(P0D50),
				.a4(P0D60),
				.a5(P0D70),
				.a6(P0E50),
				.a7(P0E60),
				.a8(P0E70),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00C50)
);

ninexnine_unit ninexnine_unit_520(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C51),
				.a1(P0C61),
				.a2(P0C71),
				.a3(P0D51),
				.a4(P0D61),
				.a5(P0D71),
				.a6(P0E51),
				.a7(P0E61),
				.a8(P0E71),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01C50)
);

ninexnine_unit ninexnine_unit_521(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C52),
				.a1(P0C62),
				.a2(P0C72),
				.a3(P0D52),
				.a4(P0D62),
				.a5(P0D72),
				.a6(P0E52),
				.a7(P0E62),
				.a8(P0E72),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02C50)
);

assign C0C50=c00C50+c01C50+c02C50;
assign A0C50=(C0C50>=0)?1:0;

ninexnine_unit ninexnine_unit_522(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C60),
				.a1(P0C70),
				.a2(P0C80),
				.a3(P0D60),
				.a4(P0D70),
				.a5(P0D80),
				.a6(P0E60),
				.a7(P0E70),
				.a8(P0E80),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00C60)
);

ninexnine_unit ninexnine_unit_523(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C61),
				.a1(P0C71),
				.a2(P0C81),
				.a3(P0D61),
				.a4(P0D71),
				.a5(P0D81),
				.a6(P0E61),
				.a7(P0E71),
				.a8(P0E81),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01C60)
);

ninexnine_unit ninexnine_unit_524(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C62),
				.a1(P0C72),
				.a2(P0C82),
				.a3(P0D62),
				.a4(P0D72),
				.a5(P0D82),
				.a6(P0E62),
				.a7(P0E72),
				.a8(P0E82),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02C60)
);

assign C0C60=c00C60+c01C60+c02C60;
assign A0C60=(C0C60>=0)?1:0;

ninexnine_unit ninexnine_unit_525(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C70),
				.a1(P0C80),
				.a2(P0C90),
				.a3(P0D70),
				.a4(P0D80),
				.a5(P0D90),
				.a6(P0E70),
				.a7(P0E80),
				.a8(P0E90),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00C70)
);

ninexnine_unit ninexnine_unit_526(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C71),
				.a1(P0C81),
				.a2(P0C91),
				.a3(P0D71),
				.a4(P0D81),
				.a5(P0D91),
				.a6(P0E71),
				.a7(P0E81),
				.a8(P0E91),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01C70)
);

ninexnine_unit ninexnine_unit_527(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C72),
				.a1(P0C82),
				.a2(P0C92),
				.a3(P0D72),
				.a4(P0D82),
				.a5(P0D92),
				.a6(P0E72),
				.a7(P0E82),
				.a8(P0E92),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02C70)
);

assign C0C70=c00C70+c01C70+c02C70;
assign A0C70=(C0C70>=0)?1:0;

ninexnine_unit ninexnine_unit_528(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C80),
				.a1(P0C90),
				.a2(P0CA0),
				.a3(P0D80),
				.a4(P0D90),
				.a5(P0DA0),
				.a6(P0E80),
				.a7(P0E90),
				.a8(P0EA0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00C80)
);

ninexnine_unit ninexnine_unit_529(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C81),
				.a1(P0C91),
				.a2(P0CA1),
				.a3(P0D81),
				.a4(P0D91),
				.a5(P0DA1),
				.a6(P0E81),
				.a7(P0E91),
				.a8(P0EA1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01C80)
);

ninexnine_unit ninexnine_unit_530(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C82),
				.a1(P0C92),
				.a2(P0CA2),
				.a3(P0D82),
				.a4(P0D92),
				.a5(P0DA2),
				.a6(P0E82),
				.a7(P0E92),
				.a8(P0EA2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02C80)
);

assign C0C80=c00C80+c01C80+c02C80;
assign A0C80=(C0C80>=0)?1:0;

ninexnine_unit ninexnine_unit_531(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C90),
				.a1(P0CA0),
				.a2(P0CB0),
				.a3(P0D90),
				.a4(P0DA0),
				.a5(P0DB0),
				.a6(P0E90),
				.a7(P0EA0),
				.a8(P0EB0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00C90)
);

ninexnine_unit ninexnine_unit_532(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C91),
				.a1(P0CA1),
				.a2(P0CB1),
				.a3(P0D91),
				.a4(P0DA1),
				.a5(P0DB1),
				.a6(P0E91),
				.a7(P0EA1),
				.a8(P0EB1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01C90)
);

ninexnine_unit ninexnine_unit_533(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C92),
				.a1(P0CA2),
				.a2(P0CB2),
				.a3(P0D92),
				.a4(P0DA2),
				.a5(P0DB2),
				.a6(P0E92),
				.a7(P0EA2),
				.a8(P0EB2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02C90)
);

assign C0C90=c00C90+c01C90+c02C90;
assign A0C90=(C0C90>=0)?1:0;

ninexnine_unit ninexnine_unit_534(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CA0),
				.a1(P0CB0),
				.a2(P0CC0),
				.a3(P0DA0),
				.a4(P0DB0),
				.a5(P0DC0),
				.a6(P0EA0),
				.a7(P0EB0),
				.a8(P0EC0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00CA0)
);

ninexnine_unit ninexnine_unit_535(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CA1),
				.a1(P0CB1),
				.a2(P0CC1),
				.a3(P0DA1),
				.a4(P0DB1),
				.a5(P0DC1),
				.a6(P0EA1),
				.a7(P0EB1),
				.a8(P0EC1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01CA0)
);

ninexnine_unit ninexnine_unit_536(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CA2),
				.a1(P0CB2),
				.a2(P0CC2),
				.a3(P0DA2),
				.a4(P0DB2),
				.a5(P0DC2),
				.a6(P0EA2),
				.a7(P0EB2),
				.a8(P0EC2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02CA0)
);

assign C0CA0=c00CA0+c01CA0+c02CA0;
assign A0CA0=(C0CA0>=0)?1:0;

ninexnine_unit ninexnine_unit_537(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CB0),
				.a1(P0CC0),
				.a2(P0CD0),
				.a3(P0DB0),
				.a4(P0DC0),
				.a5(P0DD0),
				.a6(P0EB0),
				.a7(P0EC0),
				.a8(P0ED0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00CB0)
);

ninexnine_unit ninexnine_unit_538(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CB1),
				.a1(P0CC1),
				.a2(P0CD1),
				.a3(P0DB1),
				.a4(P0DC1),
				.a5(P0DD1),
				.a6(P0EB1),
				.a7(P0EC1),
				.a8(P0ED1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01CB0)
);

ninexnine_unit ninexnine_unit_539(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CB2),
				.a1(P0CC2),
				.a2(P0CD2),
				.a3(P0DB2),
				.a4(P0DC2),
				.a5(P0DD2),
				.a6(P0EB2),
				.a7(P0EC2),
				.a8(P0ED2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02CB0)
);

assign C0CB0=c00CB0+c01CB0+c02CB0;
assign A0CB0=(C0CB0>=0)?1:0;

ninexnine_unit ninexnine_unit_540(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CC0),
				.a1(P0CD0),
				.a2(P0CE0),
				.a3(P0DC0),
				.a4(P0DD0),
				.a5(P0DE0),
				.a6(P0EC0),
				.a7(P0ED0),
				.a8(P0EE0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00CC0)
);

ninexnine_unit ninexnine_unit_541(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CC1),
				.a1(P0CD1),
				.a2(P0CE1),
				.a3(P0DC1),
				.a4(P0DD1),
				.a5(P0DE1),
				.a6(P0EC1),
				.a7(P0ED1),
				.a8(P0EE1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01CC0)
);

ninexnine_unit ninexnine_unit_542(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CC2),
				.a1(P0CD2),
				.a2(P0CE2),
				.a3(P0DC2),
				.a4(P0DD2),
				.a5(P0DE2),
				.a6(P0EC2),
				.a7(P0ED2),
				.a8(P0EE2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02CC0)
);

assign C0CC0=c00CC0+c01CC0+c02CC0;
assign A0CC0=(C0CC0>=0)?1:0;

ninexnine_unit ninexnine_unit_543(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CD0),
				.a1(P0CE0),
				.a2(P0CF0),
				.a3(P0DD0),
				.a4(P0DE0),
				.a5(P0DF0),
				.a6(P0ED0),
				.a7(P0EE0),
				.a8(P0EF0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00CD0)
);

ninexnine_unit ninexnine_unit_544(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CD1),
				.a1(P0CE1),
				.a2(P0CF1),
				.a3(P0DD1),
				.a4(P0DE1),
				.a5(P0DF1),
				.a6(P0ED1),
				.a7(P0EE1),
				.a8(P0EF1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01CD0)
);

ninexnine_unit ninexnine_unit_545(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CD2),
				.a1(P0CE2),
				.a2(P0CF2),
				.a3(P0DD2),
				.a4(P0DE2),
				.a5(P0DF2),
				.a6(P0ED2),
				.a7(P0EE2),
				.a8(P0EF2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02CD0)
);

assign C0CD0=c00CD0+c01CD0+c02CD0;
assign A0CD0=(C0CD0>=0)?1:0;

ninexnine_unit ninexnine_unit_546(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D00),
				.a1(P0D10),
				.a2(P0D20),
				.a3(P0E00),
				.a4(P0E10),
				.a5(P0E20),
				.a6(P0F00),
				.a7(P0F10),
				.a8(P0F20),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00D00)
);

ninexnine_unit ninexnine_unit_547(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D01),
				.a1(P0D11),
				.a2(P0D21),
				.a3(P0E01),
				.a4(P0E11),
				.a5(P0E21),
				.a6(P0F01),
				.a7(P0F11),
				.a8(P0F21),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01D00)
);

ninexnine_unit ninexnine_unit_548(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D02),
				.a1(P0D12),
				.a2(P0D22),
				.a3(P0E02),
				.a4(P0E12),
				.a5(P0E22),
				.a6(P0F02),
				.a7(P0F12),
				.a8(P0F22),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02D00)
);

assign C0D00=c00D00+c01D00+c02D00;
assign A0D00=(C0D00>=0)?1:0;

ninexnine_unit ninexnine_unit_549(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D10),
				.a1(P0D20),
				.a2(P0D30),
				.a3(P0E10),
				.a4(P0E20),
				.a5(P0E30),
				.a6(P0F10),
				.a7(P0F20),
				.a8(P0F30),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00D10)
);

ninexnine_unit ninexnine_unit_550(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D11),
				.a1(P0D21),
				.a2(P0D31),
				.a3(P0E11),
				.a4(P0E21),
				.a5(P0E31),
				.a6(P0F11),
				.a7(P0F21),
				.a8(P0F31),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01D10)
);

ninexnine_unit ninexnine_unit_551(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D12),
				.a1(P0D22),
				.a2(P0D32),
				.a3(P0E12),
				.a4(P0E22),
				.a5(P0E32),
				.a6(P0F12),
				.a7(P0F22),
				.a8(P0F32),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02D10)
);

assign C0D10=c00D10+c01D10+c02D10;
assign A0D10=(C0D10>=0)?1:0;

ninexnine_unit ninexnine_unit_552(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D20),
				.a1(P0D30),
				.a2(P0D40),
				.a3(P0E20),
				.a4(P0E30),
				.a5(P0E40),
				.a6(P0F20),
				.a7(P0F30),
				.a8(P0F40),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00D20)
);

ninexnine_unit ninexnine_unit_553(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D21),
				.a1(P0D31),
				.a2(P0D41),
				.a3(P0E21),
				.a4(P0E31),
				.a5(P0E41),
				.a6(P0F21),
				.a7(P0F31),
				.a8(P0F41),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01D20)
);

ninexnine_unit ninexnine_unit_554(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D22),
				.a1(P0D32),
				.a2(P0D42),
				.a3(P0E22),
				.a4(P0E32),
				.a5(P0E42),
				.a6(P0F22),
				.a7(P0F32),
				.a8(P0F42),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02D20)
);

assign C0D20=c00D20+c01D20+c02D20;
assign A0D20=(C0D20>=0)?1:0;

ninexnine_unit ninexnine_unit_555(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D30),
				.a1(P0D40),
				.a2(P0D50),
				.a3(P0E30),
				.a4(P0E40),
				.a5(P0E50),
				.a6(P0F30),
				.a7(P0F40),
				.a8(P0F50),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00D30)
);

ninexnine_unit ninexnine_unit_556(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D31),
				.a1(P0D41),
				.a2(P0D51),
				.a3(P0E31),
				.a4(P0E41),
				.a5(P0E51),
				.a6(P0F31),
				.a7(P0F41),
				.a8(P0F51),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01D30)
);

ninexnine_unit ninexnine_unit_557(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D32),
				.a1(P0D42),
				.a2(P0D52),
				.a3(P0E32),
				.a4(P0E42),
				.a5(P0E52),
				.a6(P0F32),
				.a7(P0F42),
				.a8(P0F52),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02D30)
);

assign C0D30=c00D30+c01D30+c02D30;
assign A0D30=(C0D30>=0)?1:0;

ninexnine_unit ninexnine_unit_558(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D40),
				.a1(P0D50),
				.a2(P0D60),
				.a3(P0E40),
				.a4(P0E50),
				.a5(P0E60),
				.a6(P0F40),
				.a7(P0F50),
				.a8(P0F60),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00D40)
);

ninexnine_unit ninexnine_unit_559(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D41),
				.a1(P0D51),
				.a2(P0D61),
				.a3(P0E41),
				.a4(P0E51),
				.a5(P0E61),
				.a6(P0F41),
				.a7(P0F51),
				.a8(P0F61),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01D40)
);

ninexnine_unit ninexnine_unit_560(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D42),
				.a1(P0D52),
				.a2(P0D62),
				.a3(P0E42),
				.a4(P0E52),
				.a5(P0E62),
				.a6(P0F42),
				.a7(P0F52),
				.a8(P0F62),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02D40)
);

assign C0D40=c00D40+c01D40+c02D40;
assign A0D40=(C0D40>=0)?1:0;

ninexnine_unit ninexnine_unit_561(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D50),
				.a1(P0D60),
				.a2(P0D70),
				.a3(P0E50),
				.a4(P0E60),
				.a5(P0E70),
				.a6(P0F50),
				.a7(P0F60),
				.a8(P0F70),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00D50)
);

ninexnine_unit ninexnine_unit_562(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D51),
				.a1(P0D61),
				.a2(P0D71),
				.a3(P0E51),
				.a4(P0E61),
				.a5(P0E71),
				.a6(P0F51),
				.a7(P0F61),
				.a8(P0F71),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01D50)
);

ninexnine_unit ninexnine_unit_563(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D52),
				.a1(P0D62),
				.a2(P0D72),
				.a3(P0E52),
				.a4(P0E62),
				.a5(P0E72),
				.a6(P0F52),
				.a7(P0F62),
				.a8(P0F72),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02D50)
);

assign C0D50=c00D50+c01D50+c02D50;
assign A0D50=(C0D50>=0)?1:0;

ninexnine_unit ninexnine_unit_564(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D60),
				.a1(P0D70),
				.a2(P0D80),
				.a3(P0E60),
				.a4(P0E70),
				.a5(P0E80),
				.a6(P0F60),
				.a7(P0F70),
				.a8(P0F80),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00D60)
);

ninexnine_unit ninexnine_unit_565(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D61),
				.a1(P0D71),
				.a2(P0D81),
				.a3(P0E61),
				.a4(P0E71),
				.a5(P0E81),
				.a6(P0F61),
				.a7(P0F71),
				.a8(P0F81),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01D60)
);

ninexnine_unit ninexnine_unit_566(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D62),
				.a1(P0D72),
				.a2(P0D82),
				.a3(P0E62),
				.a4(P0E72),
				.a5(P0E82),
				.a6(P0F62),
				.a7(P0F72),
				.a8(P0F82),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02D60)
);

assign C0D60=c00D60+c01D60+c02D60;
assign A0D60=(C0D60>=0)?1:0;

ninexnine_unit ninexnine_unit_567(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D70),
				.a1(P0D80),
				.a2(P0D90),
				.a3(P0E70),
				.a4(P0E80),
				.a5(P0E90),
				.a6(P0F70),
				.a7(P0F80),
				.a8(P0F90),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00D70)
);

ninexnine_unit ninexnine_unit_568(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D71),
				.a1(P0D81),
				.a2(P0D91),
				.a3(P0E71),
				.a4(P0E81),
				.a5(P0E91),
				.a6(P0F71),
				.a7(P0F81),
				.a8(P0F91),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01D70)
);

ninexnine_unit ninexnine_unit_569(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D72),
				.a1(P0D82),
				.a2(P0D92),
				.a3(P0E72),
				.a4(P0E82),
				.a5(P0E92),
				.a6(P0F72),
				.a7(P0F82),
				.a8(P0F92),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02D70)
);

assign C0D70=c00D70+c01D70+c02D70;
assign A0D70=(C0D70>=0)?1:0;

ninexnine_unit ninexnine_unit_570(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D80),
				.a1(P0D90),
				.a2(P0DA0),
				.a3(P0E80),
				.a4(P0E90),
				.a5(P0EA0),
				.a6(P0F80),
				.a7(P0F90),
				.a8(P0FA0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00D80)
);

ninexnine_unit ninexnine_unit_571(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D81),
				.a1(P0D91),
				.a2(P0DA1),
				.a3(P0E81),
				.a4(P0E91),
				.a5(P0EA1),
				.a6(P0F81),
				.a7(P0F91),
				.a8(P0FA1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01D80)
);

ninexnine_unit ninexnine_unit_572(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D82),
				.a1(P0D92),
				.a2(P0DA2),
				.a3(P0E82),
				.a4(P0E92),
				.a5(P0EA2),
				.a6(P0F82),
				.a7(P0F92),
				.a8(P0FA2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02D80)
);

assign C0D80=c00D80+c01D80+c02D80;
assign A0D80=(C0D80>=0)?1:0;

ninexnine_unit ninexnine_unit_573(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D90),
				.a1(P0DA0),
				.a2(P0DB0),
				.a3(P0E90),
				.a4(P0EA0),
				.a5(P0EB0),
				.a6(P0F90),
				.a7(P0FA0),
				.a8(P0FB0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00D90)
);

ninexnine_unit ninexnine_unit_574(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D91),
				.a1(P0DA1),
				.a2(P0DB1),
				.a3(P0E91),
				.a4(P0EA1),
				.a5(P0EB1),
				.a6(P0F91),
				.a7(P0FA1),
				.a8(P0FB1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01D90)
);

ninexnine_unit ninexnine_unit_575(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D92),
				.a1(P0DA2),
				.a2(P0DB2),
				.a3(P0E92),
				.a4(P0EA2),
				.a5(P0EB2),
				.a6(P0F92),
				.a7(P0FA2),
				.a8(P0FB2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02D90)
);

assign C0D90=c00D90+c01D90+c02D90;
assign A0D90=(C0D90>=0)?1:0;

ninexnine_unit ninexnine_unit_576(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DA0),
				.a1(P0DB0),
				.a2(P0DC0),
				.a3(P0EA0),
				.a4(P0EB0),
				.a5(P0EC0),
				.a6(P0FA0),
				.a7(P0FB0),
				.a8(P0FC0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00DA0)
);

ninexnine_unit ninexnine_unit_577(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DA1),
				.a1(P0DB1),
				.a2(P0DC1),
				.a3(P0EA1),
				.a4(P0EB1),
				.a5(P0EC1),
				.a6(P0FA1),
				.a7(P0FB1),
				.a8(P0FC1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01DA0)
);

ninexnine_unit ninexnine_unit_578(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DA2),
				.a1(P0DB2),
				.a2(P0DC2),
				.a3(P0EA2),
				.a4(P0EB2),
				.a5(P0EC2),
				.a6(P0FA2),
				.a7(P0FB2),
				.a8(P0FC2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02DA0)
);

assign C0DA0=c00DA0+c01DA0+c02DA0;
assign A0DA0=(C0DA0>=0)?1:0;

ninexnine_unit ninexnine_unit_579(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DB0),
				.a1(P0DC0),
				.a2(P0DD0),
				.a3(P0EB0),
				.a4(P0EC0),
				.a5(P0ED0),
				.a6(P0FB0),
				.a7(P0FC0),
				.a8(P0FD0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00DB0)
);

ninexnine_unit ninexnine_unit_580(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DB1),
				.a1(P0DC1),
				.a2(P0DD1),
				.a3(P0EB1),
				.a4(P0EC1),
				.a5(P0ED1),
				.a6(P0FB1),
				.a7(P0FC1),
				.a8(P0FD1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01DB0)
);

ninexnine_unit ninexnine_unit_581(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DB2),
				.a1(P0DC2),
				.a2(P0DD2),
				.a3(P0EB2),
				.a4(P0EC2),
				.a5(P0ED2),
				.a6(P0FB2),
				.a7(P0FC2),
				.a8(P0FD2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02DB0)
);

assign C0DB0=c00DB0+c01DB0+c02DB0;
assign A0DB0=(C0DB0>=0)?1:0;

ninexnine_unit ninexnine_unit_582(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DC0),
				.a1(P0DD0),
				.a2(P0DE0),
				.a3(P0EC0),
				.a4(P0ED0),
				.a5(P0EE0),
				.a6(P0FC0),
				.a7(P0FD0),
				.a8(P0FE0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00DC0)
);

ninexnine_unit ninexnine_unit_583(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DC1),
				.a1(P0DD1),
				.a2(P0DE1),
				.a3(P0EC1),
				.a4(P0ED1),
				.a5(P0EE1),
				.a6(P0FC1),
				.a7(P0FD1),
				.a8(P0FE1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01DC0)
);

ninexnine_unit ninexnine_unit_584(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DC2),
				.a1(P0DD2),
				.a2(P0DE2),
				.a3(P0EC2),
				.a4(P0ED2),
				.a5(P0EE2),
				.a6(P0FC2),
				.a7(P0FD2),
				.a8(P0FE2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02DC0)
);

assign C0DC0=c00DC0+c01DC0+c02DC0;
assign A0DC0=(C0DC0>=0)?1:0;

ninexnine_unit ninexnine_unit_585(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DD0),
				.a1(P0DE0),
				.a2(P0DF0),
				.a3(P0ED0),
				.a4(P0EE0),
				.a5(P0EF0),
				.a6(P0FD0),
				.a7(P0FE0),
				.a8(P0FF0),
				.b0(W00000),
				.b1(W00010),
				.b2(W00020),
				.b3(W00100),
				.b4(W00110),
				.b5(W00120),
				.b6(W00200),
				.b7(W00210),
				.b8(W00220),
				.c(c00DD0)
);

ninexnine_unit ninexnine_unit_586(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DD1),
				.a1(P0DE1),
				.a2(P0DF1),
				.a3(P0ED1),
				.a4(P0EE1),
				.a5(P0EF1),
				.a6(P0FD1),
				.a7(P0FE1),
				.a8(P0FF1),
				.b0(W00001),
				.b1(W00011),
				.b2(W00021),
				.b3(W00101),
				.b4(W00111),
				.b5(W00121),
				.b6(W00201),
				.b7(W00211),
				.b8(W00221),
				.c(c01DD0)
);

ninexnine_unit ninexnine_unit_587(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DD2),
				.a1(P0DE2),
				.a2(P0DF2),
				.a3(P0ED2),
				.a4(P0EE2),
				.a5(P0EF2),
				.a6(P0FD2),
				.a7(P0FE2),
				.a8(P0FF2),
				.b0(W00002),
				.b1(W00012),
				.b2(W00022),
				.b3(W00102),
				.b4(W00112),
				.b5(W00122),
				.b6(W00202),
				.b7(W00212),
				.b8(W00222),
				.c(c02DD0)
);

assign C0DD0=c00DD0+c01DD0+c02DD0;
assign A0DD0=(C0DD0>=0)?1:0;

ninexnine_unit ninexnine_unit_588(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00001)
);

ninexnine_unit ninexnine_unit_589(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01001)
);

ninexnine_unit ninexnine_unit_590(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02001)
);

assign C0001=c00001+c01001+c02001;
assign A0001=(C0001>=0)?1:0;

ninexnine_unit ninexnine_unit_591(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00011)
);

ninexnine_unit ninexnine_unit_592(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01011)
);

ninexnine_unit ninexnine_unit_593(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02011)
);

assign C0011=c00011+c01011+c02011;
assign A0011=(C0011>=0)?1:0;

ninexnine_unit ninexnine_unit_594(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00021)
);

ninexnine_unit ninexnine_unit_595(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01021)
);

ninexnine_unit ninexnine_unit_596(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02021)
);

assign C0021=c00021+c01021+c02021;
assign A0021=(C0021>=0)?1:0;

ninexnine_unit ninexnine_unit_597(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00031)
);

ninexnine_unit ninexnine_unit_598(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01031)
);

ninexnine_unit ninexnine_unit_599(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02031)
);

assign C0031=c00031+c01031+c02031;
assign A0031=(C0031>=0)?1:0;

ninexnine_unit ninexnine_unit_600(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00041)
);

ninexnine_unit ninexnine_unit_601(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01041)
);

ninexnine_unit ninexnine_unit_602(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02041)
);

assign C0041=c00041+c01041+c02041;
assign A0041=(C0041>=0)?1:0;

ninexnine_unit ninexnine_unit_603(
				.clk(clk),
				.rstn(rstn),
				.a0(P0050),
				.a1(P0060),
				.a2(P0070),
				.a3(P0150),
				.a4(P0160),
				.a5(P0170),
				.a6(P0250),
				.a7(P0260),
				.a8(P0270),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00051)
);

ninexnine_unit ninexnine_unit_604(
				.clk(clk),
				.rstn(rstn),
				.a0(P0051),
				.a1(P0061),
				.a2(P0071),
				.a3(P0151),
				.a4(P0161),
				.a5(P0171),
				.a6(P0251),
				.a7(P0261),
				.a8(P0271),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01051)
);

ninexnine_unit ninexnine_unit_605(
				.clk(clk),
				.rstn(rstn),
				.a0(P0052),
				.a1(P0062),
				.a2(P0072),
				.a3(P0152),
				.a4(P0162),
				.a5(P0172),
				.a6(P0252),
				.a7(P0262),
				.a8(P0272),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02051)
);

assign C0051=c00051+c01051+c02051;
assign A0051=(C0051>=0)?1:0;

ninexnine_unit ninexnine_unit_606(
				.clk(clk),
				.rstn(rstn),
				.a0(P0060),
				.a1(P0070),
				.a2(P0080),
				.a3(P0160),
				.a4(P0170),
				.a5(P0180),
				.a6(P0260),
				.a7(P0270),
				.a8(P0280),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00061)
);

ninexnine_unit ninexnine_unit_607(
				.clk(clk),
				.rstn(rstn),
				.a0(P0061),
				.a1(P0071),
				.a2(P0081),
				.a3(P0161),
				.a4(P0171),
				.a5(P0181),
				.a6(P0261),
				.a7(P0271),
				.a8(P0281),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01061)
);

ninexnine_unit ninexnine_unit_608(
				.clk(clk),
				.rstn(rstn),
				.a0(P0062),
				.a1(P0072),
				.a2(P0082),
				.a3(P0162),
				.a4(P0172),
				.a5(P0182),
				.a6(P0262),
				.a7(P0272),
				.a8(P0282),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02061)
);

assign C0061=c00061+c01061+c02061;
assign A0061=(C0061>=0)?1:0;

ninexnine_unit ninexnine_unit_609(
				.clk(clk),
				.rstn(rstn),
				.a0(P0070),
				.a1(P0080),
				.a2(P0090),
				.a3(P0170),
				.a4(P0180),
				.a5(P0190),
				.a6(P0270),
				.a7(P0280),
				.a8(P0290),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00071)
);

ninexnine_unit ninexnine_unit_610(
				.clk(clk),
				.rstn(rstn),
				.a0(P0071),
				.a1(P0081),
				.a2(P0091),
				.a3(P0171),
				.a4(P0181),
				.a5(P0191),
				.a6(P0271),
				.a7(P0281),
				.a8(P0291),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01071)
);

ninexnine_unit ninexnine_unit_611(
				.clk(clk),
				.rstn(rstn),
				.a0(P0072),
				.a1(P0082),
				.a2(P0092),
				.a3(P0172),
				.a4(P0182),
				.a5(P0192),
				.a6(P0272),
				.a7(P0282),
				.a8(P0292),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02071)
);

assign C0071=c00071+c01071+c02071;
assign A0071=(C0071>=0)?1:0;

ninexnine_unit ninexnine_unit_612(
				.clk(clk),
				.rstn(rstn),
				.a0(P0080),
				.a1(P0090),
				.a2(P00A0),
				.a3(P0180),
				.a4(P0190),
				.a5(P01A0),
				.a6(P0280),
				.a7(P0290),
				.a8(P02A0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00081)
);

ninexnine_unit ninexnine_unit_613(
				.clk(clk),
				.rstn(rstn),
				.a0(P0081),
				.a1(P0091),
				.a2(P00A1),
				.a3(P0181),
				.a4(P0191),
				.a5(P01A1),
				.a6(P0281),
				.a7(P0291),
				.a8(P02A1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01081)
);

ninexnine_unit ninexnine_unit_614(
				.clk(clk),
				.rstn(rstn),
				.a0(P0082),
				.a1(P0092),
				.a2(P00A2),
				.a3(P0182),
				.a4(P0192),
				.a5(P01A2),
				.a6(P0282),
				.a7(P0292),
				.a8(P02A2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02081)
);

assign C0081=c00081+c01081+c02081;
assign A0081=(C0081>=0)?1:0;

ninexnine_unit ninexnine_unit_615(
				.clk(clk),
				.rstn(rstn),
				.a0(P0090),
				.a1(P00A0),
				.a2(P00B0),
				.a3(P0190),
				.a4(P01A0),
				.a5(P01B0),
				.a6(P0290),
				.a7(P02A0),
				.a8(P02B0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00091)
);

ninexnine_unit ninexnine_unit_616(
				.clk(clk),
				.rstn(rstn),
				.a0(P0091),
				.a1(P00A1),
				.a2(P00B1),
				.a3(P0191),
				.a4(P01A1),
				.a5(P01B1),
				.a6(P0291),
				.a7(P02A1),
				.a8(P02B1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01091)
);

ninexnine_unit ninexnine_unit_617(
				.clk(clk),
				.rstn(rstn),
				.a0(P0092),
				.a1(P00A2),
				.a2(P00B2),
				.a3(P0192),
				.a4(P01A2),
				.a5(P01B2),
				.a6(P0292),
				.a7(P02A2),
				.a8(P02B2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02091)
);

assign C0091=c00091+c01091+c02091;
assign A0091=(C0091>=0)?1:0;

ninexnine_unit ninexnine_unit_618(
				.clk(clk),
				.rstn(rstn),
				.a0(P00A0),
				.a1(P00B0),
				.a2(P00C0),
				.a3(P01A0),
				.a4(P01B0),
				.a5(P01C0),
				.a6(P02A0),
				.a7(P02B0),
				.a8(P02C0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c000A1)
);

ninexnine_unit ninexnine_unit_619(
				.clk(clk),
				.rstn(rstn),
				.a0(P00A1),
				.a1(P00B1),
				.a2(P00C1),
				.a3(P01A1),
				.a4(P01B1),
				.a5(P01C1),
				.a6(P02A1),
				.a7(P02B1),
				.a8(P02C1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c010A1)
);

ninexnine_unit ninexnine_unit_620(
				.clk(clk),
				.rstn(rstn),
				.a0(P00A2),
				.a1(P00B2),
				.a2(P00C2),
				.a3(P01A2),
				.a4(P01B2),
				.a5(P01C2),
				.a6(P02A2),
				.a7(P02B2),
				.a8(P02C2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c020A1)
);

assign C00A1=c000A1+c010A1+c020A1;
assign A00A1=(C00A1>=0)?1:0;

ninexnine_unit ninexnine_unit_621(
				.clk(clk),
				.rstn(rstn),
				.a0(P00B0),
				.a1(P00C0),
				.a2(P00D0),
				.a3(P01B0),
				.a4(P01C0),
				.a5(P01D0),
				.a6(P02B0),
				.a7(P02C0),
				.a8(P02D0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c000B1)
);

ninexnine_unit ninexnine_unit_622(
				.clk(clk),
				.rstn(rstn),
				.a0(P00B1),
				.a1(P00C1),
				.a2(P00D1),
				.a3(P01B1),
				.a4(P01C1),
				.a5(P01D1),
				.a6(P02B1),
				.a7(P02C1),
				.a8(P02D1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c010B1)
);

ninexnine_unit ninexnine_unit_623(
				.clk(clk),
				.rstn(rstn),
				.a0(P00B2),
				.a1(P00C2),
				.a2(P00D2),
				.a3(P01B2),
				.a4(P01C2),
				.a5(P01D2),
				.a6(P02B2),
				.a7(P02C2),
				.a8(P02D2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c020B1)
);

assign C00B1=c000B1+c010B1+c020B1;
assign A00B1=(C00B1>=0)?1:0;

ninexnine_unit ninexnine_unit_624(
				.clk(clk),
				.rstn(rstn),
				.a0(P00C0),
				.a1(P00D0),
				.a2(P00E0),
				.a3(P01C0),
				.a4(P01D0),
				.a5(P01E0),
				.a6(P02C0),
				.a7(P02D0),
				.a8(P02E0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c000C1)
);

ninexnine_unit ninexnine_unit_625(
				.clk(clk),
				.rstn(rstn),
				.a0(P00C1),
				.a1(P00D1),
				.a2(P00E1),
				.a3(P01C1),
				.a4(P01D1),
				.a5(P01E1),
				.a6(P02C1),
				.a7(P02D1),
				.a8(P02E1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c010C1)
);

ninexnine_unit ninexnine_unit_626(
				.clk(clk),
				.rstn(rstn),
				.a0(P00C2),
				.a1(P00D2),
				.a2(P00E2),
				.a3(P01C2),
				.a4(P01D2),
				.a5(P01E2),
				.a6(P02C2),
				.a7(P02D2),
				.a8(P02E2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c020C1)
);

assign C00C1=c000C1+c010C1+c020C1;
assign A00C1=(C00C1>=0)?1:0;

ninexnine_unit ninexnine_unit_627(
				.clk(clk),
				.rstn(rstn),
				.a0(P00D0),
				.a1(P00E0),
				.a2(P00F0),
				.a3(P01D0),
				.a4(P01E0),
				.a5(P01F0),
				.a6(P02D0),
				.a7(P02E0),
				.a8(P02F0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c000D1)
);

ninexnine_unit ninexnine_unit_628(
				.clk(clk),
				.rstn(rstn),
				.a0(P00D1),
				.a1(P00E1),
				.a2(P00F1),
				.a3(P01D1),
				.a4(P01E1),
				.a5(P01F1),
				.a6(P02D1),
				.a7(P02E1),
				.a8(P02F1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c010D1)
);

ninexnine_unit ninexnine_unit_629(
				.clk(clk),
				.rstn(rstn),
				.a0(P00D2),
				.a1(P00E2),
				.a2(P00F2),
				.a3(P01D2),
				.a4(P01E2),
				.a5(P01F2),
				.a6(P02D2),
				.a7(P02E2),
				.a8(P02F2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c020D1)
);

assign C00D1=c000D1+c010D1+c020D1;
assign A00D1=(C00D1>=0)?1:0;

ninexnine_unit ninexnine_unit_630(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00101)
);

ninexnine_unit ninexnine_unit_631(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01101)
);

ninexnine_unit ninexnine_unit_632(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02101)
);

assign C0101=c00101+c01101+c02101;
assign A0101=(C0101>=0)?1:0;

ninexnine_unit ninexnine_unit_633(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00111)
);

ninexnine_unit ninexnine_unit_634(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01111)
);

ninexnine_unit ninexnine_unit_635(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02111)
);

assign C0111=c00111+c01111+c02111;
assign A0111=(C0111>=0)?1:0;

ninexnine_unit ninexnine_unit_636(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00121)
);

ninexnine_unit ninexnine_unit_637(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01121)
);

ninexnine_unit ninexnine_unit_638(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02121)
);

assign C0121=c00121+c01121+c02121;
assign A0121=(C0121>=0)?1:0;

ninexnine_unit ninexnine_unit_639(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00131)
);

ninexnine_unit ninexnine_unit_640(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01131)
);

ninexnine_unit ninexnine_unit_641(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02131)
);

assign C0131=c00131+c01131+c02131;
assign A0131=(C0131>=0)?1:0;

ninexnine_unit ninexnine_unit_642(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00141)
);

ninexnine_unit ninexnine_unit_643(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01141)
);

ninexnine_unit ninexnine_unit_644(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02141)
);

assign C0141=c00141+c01141+c02141;
assign A0141=(C0141>=0)?1:0;

ninexnine_unit ninexnine_unit_645(
				.clk(clk),
				.rstn(rstn),
				.a0(P0150),
				.a1(P0160),
				.a2(P0170),
				.a3(P0250),
				.a4(P0260),
				.a5(P0270),
				.a6(P0350),
				.a7(P0360),
				.a8(P0370),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00151)
);

ninexnine_unit ninexnine_unit_646(
				.clk(clk),
				.rstn(rstn),
				.a0(P0151),
				.a1(P0161),
				.a2(P0171),
				.a3(P0251),
				.a4(P0261),
				.a5(P0271),
				.a6(P0351),
				.a7(P0361),
				.a8(P0371),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01151)
);

ninexnine_unit ninexnine_unit_647(
				.clk(clk),
				.rstn(rstn),
				.a0(P0152),
				.a1(P0162),
				.a2(P0172),
				.a3(P0252),
				.a4(P0262),
				.a5(P0272),
				.a6(P0352),
				.a7(P0362),
				.a8(P0372),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02151)
);

assign C0151=c00151+c01151+c02151;
assign A0151=(C0151>=0)?1:0;

ninexnine_unit ninexnine_unit_648(
				.clk(clk),
				.rstn(rstn),
				.a0(P0160),
				.a1(P0170),
				.a2(P0180),
				.a3(P0260),
				.a4(P0270),
				.a5(P0280),
				.a6(P0360),
				.a7(P0370),
				.a8(P0380),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00161)
);

ninexnine_unit ninexnine_unit_649(
				.clk(clk),
				.rstn(rstn),
				.a0(P0161),
				.a1(P0171),
				.a2(P0181),
				.a3(P0261),
				.a4(P0271),
				.a5(P0281),
				.a6(P0361),
				.a7(P0371),
				.a8(P0381),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01161)
);

ninexnine_unit ninexnine_unit_650(
				.clk(clk),
				.rstn(rstn),
				.a0(P0162),
				.a1(P0172),
				.a2(P0182),
				.a3(P0262),
				.a4(P0272),
				.a5(P0282),
				.a6(P0362),
				.a7(P0372),
				.a8(P0382),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02161)
);

assign C0161=c00161+c01161+c02161;
assign A0161=(C0161>=0)?1:0;

ninexnine_unit ninexnine_unit_651(
				.clk(clk),
				.rstn(rstn),
				.a0(P0170),
				.a1(P0180),
				.a2(P0190),
				.a3(P0270),
				.a4(P0280),
				.a5(P0290),
				.a6(P0370),
				.a7(P0380),
				.a8(P0390),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00171)
);

ninexnine_unit ninexnine_unit_652(
				.clk(clk),
				.rstn(rstn),
				.a0(P0171),
				.a1(P0181),
				.a2(P0191),
				.a3(P0271),
				.a4(P0281),
				.a5(P0291),
				.a6(P0371),
				.a7(P0381),
				.a8(P0391),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01171)
);

ninexnine_unit ninexnine_unit_653(
				.clk(clk),
				.rstn(rstn),
				.a0(P0172),
				.a1(P0182),
				.a2(P0192),
				.a3(P0272),
				.a4(P0282),
				.a5(P0292),
				.a6(P0372),
				.a7(P0382),
				.a8(P0392),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02171)
);

assign C0171=c00171+c01171+c02171;
assign A0171=(C0171>=0)?1:0;

ninexnine_unit ninexnine_unit_654(
				.clk(clk),
				.rstn(rstn),
				.a0(P0180),
				.a1(P0190),
				.a2(P01A0),
				.a3(P0280),
				.a4(P0290),
				.a5(P02A0),
				.a6(P0380),
				.a7(P0390),
				.a8(P03A0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00181)
);

ninexnine_unit ninexnine_unit_655(
				.clk(clk),
				.rstn(rstn),
				.a0(P0181),
				.a1(P0191),
				.a2(P01A1),
				.a3(P0281),
				.a4(P0291),
				.a5(P02A1),
				.a6(P0381),
				.a7(P0391),
				.a8(P03A1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01181)
);

ninexnine_unit ninexnine_unit_656(
				.clk(clk),
				.rstn(rstn),
				.a0(P0182),
				.a1(P0192),
				.a2(P01A2),
				.a3(P0282),
				.a4(P0292),
				.a5(P02A2),
				.a6(P0382),
				.a7(P0392),
				.a8(P03A2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02181)
);

assign C0181=c00181+c01181+c02181;
assign A0181=(C0181>=0)?1:0;

ninexnine_unit ninexnine_unit_657(
				.clk(clk),
				.rstn(rstn),
				.a0(P0190),
				.a1(P01A0),
				.a2(P01B0),
				.a3(P0290),
				.a4(P02A0),
				.a5(P02B0),
				.a6(P0390),
				.a7(P03A0),
				.a8(P03B0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00191)
);

ninexnine_unit ninexnine_unit_658(
				.clk(clk),
				.rstn(rstn),
				.a0(P0191),
				.a1(P01A1),
				.a2(P01B1),
				.a3(P0291),
				.a4(P02A1),
				.a5(P02B1),
				.a6(P0391),
				.a7(P03A1),
				.a8(P03B1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01191)
);

ninexnine_unit ninexnine_unit_659(
				.clk(clk),
				.rstn(rstn),
				.a0(P0192),
				.a1(P01A2),
				.a2(P01B2),
				.a3(P0292),
				.a4(P02A2),
				.a5(P02B2),
				.a6(P0392),
				.a7(P03A2),
				.a8(P03B2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02191)
);

assign C0191=c00191+c01191+c02191;
assign A0191=(C0191>=0)?1:0;

ninexnine_unit ninexnine_unit_660(
				.clk(clk),
				.rstn(rstn),
				.a0(P01A0),
				.a1(P01B0),
				.a2(P01C0),
				.a3(P02A0),
				.a4(P02B0),
				.a5(P02C0),
				.a6(P03A0),
				.a7(P03B0),
				.a8(P03C0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c001A1)
);

ninexnine_unit ninexnine_unit_661(
				.clk(clk),
				.rstn(rstn),
				.a0(P01A1),
				.a1(P01B1),
				.a2(P01C1),
				.a3(P02A1),
				.a4(P02B1),
				.a5(P02C1),
				.a6(P03A1),
				.a7(P03B1),
				.a8(P03C1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c011A1)
);

ninexnine_unit ninexnine_unit_662(
				.clk(clk),
				.rstn(rstn),
				.a0(P01A2),
				.a1(P01B2),
				.a2(P01C2),
				.a3(P02A2),
				.a4(P02B2),
				.a5(P02C2),
				.a6(P03A2),
				.a7(P03B2),
				.a8(P03C2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c021A1)
);

assign C01A1=c001A1+c011A1+c021A1;
assign A01A1=(C01A1>=0)?1:0;

ninexnine_unit ninexnine_unit_663(
				.clk(clk),
				.rstn(rstn),
				.a0(P01B0),
				.a1(P01C0),
				.a2(P01D0),
				.a3(P02B0),
				.a4(P02C0),
				.a5(P02D0),
				.a6(P03B0),
				.a7(P03C0),
				.a8(P03D0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c001B1)
);

ninexnine_unit ninexnine_unit_664(
				.clk(clk),
				.rstn(rstn),
				.a0(P01B1),
				.a1(P01C1),
				.a2(P01D1),
				.a3(P02B1),
				.a4(P02C1),
				.a5(P02D1),
				.a6(P03B1),
				.a7(P03C1),
				.a8(P03D1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c011B1)
);

ninexnine_unit ninexnine_unit_665(
				.clk(clk),
				.rstn(rstn),
				.a0(P01B2),
				.a1(P01C2),
				.a2(P01D2),
				.a3(P02B2),
				.a4(P02C2),
				.a5(P02D2),
				.a6(P03B2),
				.a7(P03C2),
				.a8(P03D2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c021B1)
);

assign C01B1=c001B1+c011B1+c021B1;
assign A01B1=(C01B1>=0)?1:0;

ninexnine_unit ninexnine_unit_666(
				.clk(clk),
				.rstn(rstn),
				.a0(P01C0),
				.a1(P01D0),
				.a2(P01E0),
				.a3(P02C0),
				.a4(P02D0),
				.a5(P02E0),
				.a6(P03C0),
				.a7(P03D0),
				.a8(P03E0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c001C1)
);

ninexnine_unit ninexnine_unit_667(
				.clk(clk),
				.rstn(rstn),
				.a0(P01C1),
				.a1(P01D1),
				.a2(P01E1),
				.a3(P02C1),
				.a4(P02D1),
				.a5(P02E1),
				.a6(P03C1),
				.a7(P03D1),
				.a8(P03E1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c011C1)
);

ninexnine_unit ninexnine_unit_668(
				.clk(clk),
				.rstn(rstn),
				.a0(P01C2),
				.a1(P01D2),
				.a2(P01E2),
				.a3(P02C2),
				.a4(P02D2),
				.a5(P02E2),
				.a6(P03C2),
				.a7(P03D2),
				.a8(P03E2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c021C1)
);

assign C01C1=c001C1+c011C1+c021C1;
assign A01C1=(C01C1>=0)?1:0;

ninexnine_unit ninexnine_unit_669(
				.clk(clk),
				.rstn(rstn),
				.a0(P01D0),
				.a1(P01E0),
				.a2(P01F0),
				.a3(P02D0),
				.a4(P02E0),
				.a5(P02F0),
				.a6(P03D0),
				.a7(P03E0),
				.a8(P03F0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c001D1)
);

ninexnine_unit ninexnine_unit_670(
				.clk(clk),
				.rstn(rstn),
				.a0(P01D1),
				.a1(P01E1),
				.a2(P01F1),
				.a3(P02D1),
				.a4(P02E1),
				.a5(P02F1),
				.a6(P03D1),
				.a7(P03E1),
				.a8(P03F1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c011D1)
);

ninexnine_unit ninexnine_unit_671(
				.clk(clk),
				.rstn(rstn),
				.a0(P01D2),
				.a1(P01E2),
				.a2(P01F2),
				.a3(P02D2),
				.a4(P02E2),
				.a5(P02F2),
				.a6(P03D2),
				.a7(P03E2),
				.a8(P03F2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c021D1)
);

assign C01D1=c001D1+c011D1+c021D1;
assign A01D1=(C01D1>=0)?1:0;

ninexnine_unit ninexnine_unit_672(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00201)
);

ninexnine_unit ninexnine_unit_673(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01201)
);

ninexnine_unit ninexnine_unit_674(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02201)
);

assign C0201=c00201+c01201+c02201;
assign A0201=(C0201>=0)?1:0;

ninexnine_unit ninexnine_unit_675(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00211)
);

ninexnine_unit ninexnine_unit_676(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01211)
);

ninexnine_unit ninexnine_unit_677(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02211)
);

assign C0211=c00211+c01211+c02211;
assign A0211=(C0211>=0)?1:0;

ninexnine_unit ninexnine_unit_678(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00221)
);

ninexnine_unit ninexnine_unit_679(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01221)
);

ninexnine_unit ninexnine_unit_680(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02221)
);

assign C0221=c00221+c01221+c02221;
assign A0221=(C0221>=0)?1:0;

ninexnine_unit ninexnine_unit_681(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00231)
);

ninexnine_unit ninexnine_unit_682(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01231)
);

ninexnine_unit ninexnine_unit_683(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02231)
);

assign C0231=c00231+c01231+c02231;
assign A0231=(C0231>=0)?1:0;

ninexnine_unit ninexnine_unit_684(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00241)
);

ninexnine_unit ninexnine_unit_685(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01241)
);

ninexnine_unit ninexnine_unit_686(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02241)
);

assign C0241=c00241+c01241+c02241;
assign A0241=(C0241>=0)?1:0;

ninexnine_unit ninexnine_unit_687(
				.clk(clk),
				.rstn(rstn),
				.a0(P0250),
				.a1(P0260),
				.a2(P0270),
				.a3(P0350),
				.a4(P0360),
				.a5(P0370),
				.a6(P0450),
				.a7(P0460),
				.a8(P0470),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00251)
);

ninexnine_unit ninexnine_unit_688(
				.clk(clk),
				.rstn(rstn),
				.a0(P0251),
				.a1(P0261),
				.a2(P0271),
				.a3(P0351),
				.a4(P0361),
				.a5(P0371),
				.a6(P0451),
				.a7(P0461),
				.a8(P0471),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01251)
);

ninexnine_unit ninexnine_unit_689(
				.clk(clk),
				.rstn(rstn),
				.a0(P0252),
				.a1(P0262),
				.a2(P0272),
				.a3(P0352),
				.a4(P0362),
				.a5(P0372),
				.a6(P0452),
				.a7(P0462),
				.a8(P0472),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02251)
);

assign C0251=c00251+c01251+c02251;
assign A0251=(C0251>=0)?1:0;

ninexnine_unit ninexnine_unit_690(
				.clk(clk),
				.rstn(rstn),
				.a0(P0260),
				.a1(P0270),
				.a2(P0280),
				.a3(P0360),
				.a4(P0370),
				.a5(P0380),
				.a6(P0460),
				.a7(P0470),
				.a8(P0480),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00261)
);

ninexnine_unit ninexnine_unit_691(
				.clk(clk),
				.rstn(rstn),
				.a0(P0261),
				.a1(P0271),
				.a2(P0281),
				.a3(P0361),
				.a4(P0371),
				.a5(P0381),
				.a6(P0461),
				.a7(P0471),
				.a8(P0481),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01261)
);

ninexnine_unit ninexnine_unit_692(
				.clk(clk),
				.rstn(rstn),
				.a0(P0262),
				.a1(P0272),
				.a2(P0282),
				.a3(P0362),
				.a4(P0372),
				.a5(P0382),
				.a6(P0462),
				.a7(P0472),
				.a8(P0482),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02261)
);

assign C0261=c00261+c01261+c02261;
assign A0261=(C0261>=0)?1:0;

ninexnine_unit ninexnine_unit_693(
				.clk(clk),
				.rstn(rstn),
				.a0(P0270),
				.a1(P0280),
				.a2(P0290),
				.a3(P0370),
				.a4(P0380),
				.a5(P0390),
				.a6(P0470),
				.a7(P0480),
				.a8(P0490),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00271)
);

ninexnine_unit ninexnine_unit_694(
				.clk(clk),
				.rstn(rstn),
				.a0(P0271),
				.a1(P0281),
				.a2(P0291),
				.a3(P0371),
				.a4(P0381),
				.a5(P0391),
				.a6(P0471),
				.a7(P0481),
				.a8(P0491),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01271)
);

ninexnine_unit ninexnine_unit_695(
				.clk(clk),
				.rstn(rstn),
				.a0(P0272),
				.a1(P0282),
				.a2(P0292),
				.a3(P0372),
				.a4(P0382),
				.a5(P0392),
				.a6(P0472),
				.a7(P0482),
				.a8(P0492),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02271)
);

assign C0271=c00271+c01271+c02271;
assign A0271=(C0271>=0)?1:0;

ninexnine_unit ninexnine_unit_696(
				.clk(clk),
				.rstn(rstn),
				.a0(P0280),
				.a1(P0290),
				.a2(P02A0),
				.a3(P0380),
				.a4(P0390),
				.a5(P03A0),
				.a6(P0480),
				.a7(P0490),
				.a8(P04A0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00281)
);

ninexnine_unit ninexnine_unit_697(
				.clk(clk),
				.rstn(rstn),
				.a0(P0281),
				.a1(P0291),
				.a2(P02A1),
				.a3(P0381),
				.a4(P0391),
				.a5(P03A1),
				.a6(P0481),
				.a7(P0491),
				.a8(P04A1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01281)
);

ninexnine_unit ninexnine_unit_698(
				.clk(clk),
				.rstn(rstn),
				.a0(P0282),
				.a1(P0292),
				.a2(P02A2),
				.a3(P0382),
				.a4(P0392),
				.a5(P03A2),
				.a6(P0482),
				.a7(P0492),
				.a8(P04A2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02281)
);

assign C0281=c00281+c01281+c02281;
assign A0281=(C0281>=0)?1:0;

ninexnine_unit ninexnine_unit_699(
				.clk(clk),
				.rstn(rstn),
				.a0(P0290),
				.a1(P02A0),
				.a2(P02B0),
				.a3(P0390),
				.a4(P03A0),
				.a5(P03B0),
				.a6(P0490),
				.a7(P04A0),
				.a8(P04B0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00291)
);

ninexnine_unit ninexnine_unit_700(
				.clk(clk),
				.rstn(rstn),
				.a0(P0291),
				.a1(P02A1),
				.a2(P02B1),
				.a3(P0391),
				.a4(P03A1),
				.a5(P03B1),
				.a6(P0491),
				.a7(P04A1),
				.a8(P04B1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01291)
);

ninexnine_unit ninexnine_unit_701(
				.clk(clk),
				.rstn(rstn),
				.a0(P0292),
				.a1(P02A2),
				.a2(P02B2),
				.a3(P0392),
				.a4(P03A2),
				.a5(P03B2),
				.a6(P0492),
				.a7(P04A2),
				.a8(P04B2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02291)
);

assign C0291=c00291+c01291+c02291;
assign A0291=(C0291>=0)?1:0;

ninexnine_unit ninexnine_unit_702(
				.clk(clk),
				.rstn(rstn),
				.a0(P02A0),
				.a1(P02B0),
				.a2(P02C0),
				.a3(P03A0),
				.a4(P03B0),
				.a5(P03C0),
				.a6(P04A0),
				.a7(P04B0),
				.a8(P04C0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c002A1)
);

ninexnine_unit ninexnine_unit_703(
				.clk(clk),
				.rstn(rstn),
				.a0(P02A1),
				.a1(P02B1),
				.a2(P02C1),
				.a3(P03A1),
				.a4(P03B1),
				.a5(P03C1),
				.a6(P04A1),
				.a7(P04B1),
				.a8(P04C1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c012A1)
);

ninexnine_unit ninexnine_unit_704(
				.clk(clk),
				.rstn(rstn),
				.a0(P02A2),
				.a1(P02B2),
				.a2(P02C2),
				.a3(P03A2),
				.a4(P03B2),
				.a5(P03C2),
				.a6(P04A2),
				.a7(P04B2),
				.a8(P04C2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c022A1)
);

assign C02A1=c002A1+c012A1+c022A1;
assign A02A1=(C02A1>=0)?1:0;

ninexnine_unit ninexnine_unit_705(
				.clk(clk),
				.rstn(rstn),
				.a0(P02B0),
				.a1(P02C0),
				.a2(P02D0),
				.a3(P03B0),
				.a4(P03C0),
				.a5(P03D0),
				.a6(P04B0),
				.a7(P04C0),
				.a8(P04D0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c002B1)
);

ninexnine_unit ninexnine_unit_706(
				.clk(clk),
				.rstn(rstn),
				.a0(P02B1),
				.a1(P02C1),
				.a2(P02D1),
				.a3(P03B1),
				.a4(P03C1),
				.a5(P03D1),
				.a6(P04B1),
				.a7(P04C1),
				.a8(P04D1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c012B1)
);

ninexnine_unit ninexnine_unit_707(
				.clk(clk),
				.rstn(rstn),
				.a0(P02B2),
				.a1(P02C2),
				.a2(P02D2),
				.a3(P03B2),
				.a4(P03C2),
				.a5(P03D2),
				.a6(P04B2),
				.a7(P04C2),
				.a8(P04D2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c022B1)
);

assign C02B1=c002B1+c012B1+c022B1;
assign A02B1=(C02B1>=0)?1:0;

ninexnine_unit ninexnine_unit_708(
				.clk(clk),
				.rstn(rstn),
				.a0(P02C0),
				.a1(P02D0),
				.a2(P02E0),
				.a3(P03C0),
				.a4(P03D0),
				.a5(P03E0),
				.a6(P04C0),
				.a7(P04D0),
				.a8(P04E0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c002C1)
);

ninexnine_unit ninexnine_unit_709(
				.clk(clk),
				.rstn(rstn),
				.a0(P02C1),
				.a1(P02D1),
				.a2(P02E1),
				.a3(P03C1),
				.a4(P03D1),
				.a5(P03E1),
				.a6(P04C1),
				.a7(P04D1),
				.a8(P04E1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c012C1)
);

ninexnine_unit ninexnine_unit_710(
				.clk(clk),
				.rstn(rstn),
				.a0(P02C2),
				.a1(P02D2),
				.a2(P02E2),
				.a3(P03C2),
				.a4(P03D2),
				.a5(P03E2),
				.a6(P04C2),
				.a7(P04D2),
				.a8(P04E2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c022C1)
);

assign C02C1=c002C1+c012C1+c022C1;
assign A02C1=(C02C1>=0)?1:0;

ninexnine_unit ninexnine_unit_711(
				.clk(clk),
				.rstn(rstn),
				.a0(P02D0),
				.a1(P02E0),
				.a2(P02F0),
				.a3(P03D0),
				.a4(P03E0),
				.a5(P03F0),
				.a6(P04D0),
				.a7(P04E0),
				.a8(P04F0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c002D1)
);

ninexnine_unit ninexnine_unit_712(
				.clk(clk),
				.rstn(rstn),
				.a0(P02D1),
				.a1(P02E1),
				.a2(P02F1),
				.a3(P03D1),
				.a4(P03E1),
				.a5(P03F1),
				.a6(P04D1),
				.a7(P04E1),
				.a8(P04F1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c012D1)
);

ninexnine_unit ninexnine_unit_713(
				.clk(clk),
				.rstn(rstn),
				.a0(P02D2),
				.a1(P02E2),
				.a2(P02F2),
				.a3(P03D2),
				.a4(P03E2),
				.a5(P03F2),
				.a6(P04D2),
				.a7(P04E2),
				.a8(P04F2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c022D1)
);

assign C02D1=c002D1+c012D1+c022D1;
assign A02D1=(C02D1>=0)?1:0;

ninexnine_unit ninexnine_unit_714(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00301)
);

ninexnine_unit ninexnine_unit_715(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01301)
);

ninexnine_unit ninexnine_unit_716(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02301)
);

assign C0301=c00301+c01301+c02301;
assign A0301=(C0301>=0)?1:0;

ninexnine_unit ninexnine_unit_717(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00311)
);

ninexnine_unit ninexnine_unit_718(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01311)
);

ninexnine_unit ninexnine_unit_719(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02311)
);

assign C0311=c00311+c01311+c02311;
assign A0311=(C0311>=0)?1:0;

ninexnine_unit ninexnine_unit_720(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00321)
);

ninexnine_unit ninexnine_unit_721(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01321)
);

ninexnine_unit ninexnine_unit_722(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02321)
);

assign C0321=c00321+c01321+c02321;
assign A0321=(C0321>=0)?1:0;

ninexnine_unit ninexnine_unit_723(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00331)
);

ninexnine_unit ninexnine_unit_724(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01331)
);

ninexnine_unit ninexnine_unit_725(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02331)
);

assign C0331=c00331+c01331+c02331;
assign A0331=(C0331>=0)?1:0;

ninexnine_unit ninexnine_unit_726(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00341)
);

ninexnine_unit ninexnine_unit_727(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01341)
);

ninexnine_unit ninexnine_unit_728(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02341)
);

assign C0341=c00341+c01341+c02341;
assign A0341=(C0341>=0)?1:0;

ninexnine_unit ninexnine_unit_729(
				.clk(clk),
				.rstn(rstn),
				.a0(P0350),
				.a1(P0360),
				.a2(P0370),
				.a3(P0450),
				.a4(P0460),
				.a5(P0470),
				.a6(P0550),
				.a7(P0560),
				.a8(P0570),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00351)
);

ninexnine_unit ninexnine_unit_730(
				.clk(clk),
				.rstn(rstn),
				.a0(P0351),
				.a1(P0361),
				.a2(P0371),
				.a3(P0451),
				.a4(P0461),
				.a5(P0471),
				.a6(P0551),
				.a7(P0561),
				.a8(P0571),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01351)
);

ninexnine_unit ninexnine_unit_731(
				.clk(clk),
				.rstn(rstn),
				.a0(P0352),
				.a1(P0362),
				.a2(P0372),
				.a3(P0452),
				.a4(P0462),
				.a5(P0472),
				.a6(P0552),
				.a7(P0562),
				.a8(P0572),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02351)
);

assign C0351=c00351+c01351+c02351;
assign A0351=(C0351>=0)?1:0;

ninexnine_unit ninexnine_unit_732(
				.clk(clk),
				.rstn(rstn),
				.a0(P0360),
				.a1(P0370),
				.a2(P0380),
				.a3(P0460),
				.a4(P0470),
				.a5(P0480),
				.a6(P0560),
				.a7(P0570),
				.a8(P0580),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00361)
);

ninexnine_unit ninexnine_unit_733(
				.clk(clk),
				.rstn(rstn),
				.a0(P0361),
				.a1(P0371),
				.a2(P0381),
				.a3(P0461),
				.a4(P0471),
				.a5(P0481),
				.a6(P0561),
				.a7(P0571),
				.a8(P0581),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01361)
);

ninexnine_unit ninexnine_unit_734(
				.clk(clk),
				.rstn(rstn),
				.a0(P0362),
				.a1(P0372),
				.a2(P0382),
				.a3(P0462),
				.a4(P0472),
				.a5(P0482),
				.a6(P0562),
				.a7(P0572),
				.a8(P0582),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02361)
);

assign C0361=c00361+c01361+c02361;
assign A0361=(C0361>=0)?1:0;

ninexnine_unit ninexnine_unit_735(
				.clk(clk),
				.rstn(rstn),
				.a0(P0370),
				.a1(P0380),
				.a2(P0390),
				.a3(P0470),
				.a4(P0480),
				.a5(P0490),
				.a6(P0570),
				.a7(P0580),
				.a8(P0590),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00371)
);

ninexnine_unit ninexnine_unit_736(
				.clk(clk),
				.rstn(rstn),
				.a0(P0371),
				.a1(P0381),
				.a2(P0391),
				.a3(P0471),
				.a4(P0481),
				.a5(P0491),
				.a6(P0571),
				.a7(P0581),
				.a8(P0591),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01371)
);

ninexnine_unit ninexnine_unit_737(
				.clk(clk),
				.rstn(rstn),
				.a0(P0372),
				.a1(P0382),
				.a2(P0392),
				.a3(P0472),
				.a4(P0482),
				.a5(P0492),
				.a6(P0572),
				.a7(P0582),
				.a8(P0592),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02371)
);

assign C0371=c00371+c01371+c02371;
assign A0371=(C0371>=0)?1:0;

ninexnine_unit ninexnine_unit_738(
				.clk(clk),
				.rstn(rstn),
				.a0(P0380),
				.a1(P0390),
				.a2(P03A0),
				.a3(P0480),
				.a4(P0490),
				.a5(P04A0),
				.a6(P0580),
				.a7(P0590),
				.a8(P05A0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00381)
);

ninexnine_unit ninexnine_unit_739(
				.clk(clk),
				.rstn(rstn),
				.a0(P0381),
				.a1(P0391),
				.a2(P03A1),
				.a3(P0481),
				.a4(P0491),
				.a5(P04A1),
				.a6(P0581),
				.a7(P0591),
				.a8(P05A1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01381)
);

ninexnine_unit ninexnine_unit_740(
				.clk(clk),
				.rstn(rstn),
				.a0(P0382),
				.a1(P0392),
				.a2(P03A2),
				.a3(P0482),
				.a4(P0492),
				.a5(P04A2),
				.a6(P0582),
				.a7(P0592),
				.a8(P05A2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02381)
);

assign C0381=c00381+c01381+c02381;
assign A0381=(C0381>=0)?1:0;

ninexnine_unit ninexnine_unit_741(
				.clk(clk),
				.rstn(rstn),
				.a0(P0390),
				.a1(P03A0),
				.a2(P03B0),
				.a3(P0490),
				.a4(P04A0),
				.a5(P04B0),
				.a6(P0590),
				.a7(P05A0),
				.a8(P05B0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00391)
);

ninexnine_unit ninexnine_unit_742(
				.clk(clk),
				.rstn(rstn),
				.a0(P0391),
				.a1(P03A1),
				.a2(P03B1),
				.a3(P0491),
				.a4(P04A1),
				.a5(P04B1),
				.a6(P0591),
				.a7(P05A1),
				.a8(P05B1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01391)
);

ninexnine_unit ninexnine_unit_743(
				.clk(clk),
				.rstn(rstn),
				.a0(P0392),
				.a1(P03A2),
				.a2(P03B2),
				.a3(P0492),
				.a4(P04A2),
				.a5(P04B2),
				.a6(P0592),
				.a7(P05A2),
				.a8(P05B2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02391)
);

assign C0391=c00391+c01391+c02391;
assign A0391=(C0391>=0)?1:0;

ninexnine_unit ninexnine_unit_744(
				.clk(clk),
				.rstn(rstn),
				.a0(P03A0),
				.a1(P03B0),
				.a2(P03C0),
				.a3(P04A0),
				.a4(P04B0),
				.a5(P04C0),
				.a6(P05A0),
				.a7(P05B0),
				.a8(P05C0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c003A1)
);

ninexnine_unit ninexnine_unit_745(
				.clk(clk),
				.rstn(rstn),
				.a0(P03A1),
				.a1(P03B1),
				.a2(P03C1),
				.a3(P04A1),
				.a4(P04B1),
				.a5(P04C1),
				.a6(P05A1),
				.a7(P05B1),
				.a8(P05C1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c013A1)
);

ninexnine_unit ninexnine_unit_746(
				.clk(clk),
				.rstn(rstn),
				.a0(P03A2),
				.a1(P03B2),
				.a2(P03C2),
				.a3(P04A2),
				.a4(P04B2),
				.a5(P04C2),
				.a6(P05A2),
				.a7(P05B2),
				.a8(P05C2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c023A1)
);

assign C03A1=c003A1+c013A1+c023A1;
assign A03A1=(C03A1>=0)?1:0;

ninexnine_unit ninexnine_unit_747(
				.clk(clk),
				.rstn(rstn),
				.a0(P03B0),
				.a1(P03C0),
				.a2(P03D0),
				.a3(P04B0),
				.a4(P04C0),
				.a5(P04D0),
				.a6(P05B0),
				.a7(P05C0),
				.a8(P05D0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c003B1)
);

ninexnine_unit ninexnine_unit_748(
				.clk(clk),
				.rstn(rstn),
				.a0(P03B1),
				.a1(P03C1),
				.a2(P03D1),
				.a3(P04B1),
				.a4(P04C1),
				.a5(P04D1),
				.a6(P05B1),
				.a7(P05C1),
				.a8(P05D1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c013B1)
);

ninexnine_unit ninexnine_unit_749(
				.clk(clk),
				.rstn(rstn),
				.a0(P03B2),
				.a1(P03C2),
				.a2(P03D2),
				.a3(P04B2),
				.a4(P04C2),
				.a5(P04D2),
				.a6(P05B2),
				.a7(P05C2),
				.a8(P05D2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c023B1)
);

assign C03B1=c003B1+c013B1+c023B1;
assign A03B1=(C03B1>=0)?1:0;

ninexnine_unit ninexnine_unit_750(
				.clk(clk),
				.rstn(rstn),
				.a0(P03C0),
				.a1(P03D0),
				.a2(P03E0),
				.a3(P04C0),
				.a4(P04D0),
				.a5(P04E0),
				.a6(P05C0),
				.a7(P05D0),
				.a8(P05E0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c003C1)
);

ninexnine_unit ninexnine_unit_751(
				.clk(clk),
				.rstn(rstn),
				.a0(P03C1),
				.a1(P03D1),
				.a2(P03E1),
				.a3(P04C1),
				.a4(P04D1),
				.a5(P04E1),
				.a6(P05C1),
				.a7(P05D1),
				.a8(P05E1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c013C1)
);

ninexnine_unit ninexnine_unit_752(
				.clk(clk),
				.rstn(rstn),
				.a0(P03C2),
				.a1(P03D2),
				.a2(P03E2),
				.a3(P04C2),
				.a4(P04D2),
				.a5(P04E2),
				.a6(P05C2),
				.a7(P05D2),
				.a8(P05E2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c023C1)
);

assign C03C1=c003C1+c013C1+c023C1;
assign A03C1=(C03C1>=0)?1:0;

ninexnine_unit ninexnine_unit_753(
				.clk(clk),
				.rstn(rstn),
				.a0(P03D0),
				.a1(P03E0),
				.a2(P03F0),
				.a3(P04D0),
				.a4(P04E0),
				.a5(P04F0),
				.a6(P05D0),
				.a7(P05E0),
				.a8(P05F0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c003D1)
);

ninexnine_unit ninexnine_unit_754(
				.clk(clk),
				.rstn(rstn),
				.a0(P03D1),
				.a1(P03E1),
				.a2(P03F1),
				.a3(P04D1),
				.a4(P04E1),
				.a5(P04F1),
				.a6(P05D1),
				.a7(P05E1),
				.a8(P05F1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c013D1)
);

ninexnine_unit ninexnine_unit_755(
				.clk(clk),
				.rstn(rstn),
				.a0(P03D2),
				.a1(P03E2),
				.a2(P03F2),
				.a3(P04D2),
				.a4(P04E2),
				.a5(P04F2),
				.a6(P05D2),
				.a7(P05E2),
				.a8(P05F2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c023D1)
);

assign C03D1=c003D1+c013D1+c023D1;
assign A03D1=(C03D1>=0)?1:0;

ninexnine_unit ninexnine_unit_756(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00401)
);

ninexnine_unit ninexnine_unit_757(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01401)
);

ninexnine_unit ninexnine_unit_758(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02401)
);

assign C0401=c00401+c01401+c02401;
assign A0401=(C0401>=0)?1:0;

ninexnine_unit ninexnine_unit_759(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00411)
);

ninexnine_unit ninexnine_unit_760(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01411)
);

ninexnine_unit ninexnine_unit_761(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02411)
);

assign C0411=c00411+c01411+c02411;
assign A0411=(C0411>=0)?1:0;

ninexnine_unit ninexnine_unit_762(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00421)
);

ninexnine_unit ninexnine_unit_763(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01421)
);

ninexnine_unit ninexnine_unit_764(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02421)
);

assign C0421=c00421+c01421+c02421;
assign A0421=(C0421>=0)?1:0;

ninexnine_unit ninexnine_unit_765(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00431)
);

ninexnine_unit ninexnine_unit_766(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01431)
);

ninexnine_unit ninexnine_unit_767(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02431)
);

assign C0431=c00431+c01431+c02431;
assign A0431=(C0431>=0)?1:0;

ninexnine_unit ninexnine_unit_768(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00441)
);

ninexnine_unit ninexnine_unit_769(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01441)
);

ninexnine_unit ninexnine_unit_770(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02441)
);

assign C0441=c00441+c01441+c02441;
assign A0441=(C0441>=0)?1:0;

ninexnine_unit ninexnine_unit_771(
				.clk(clk),
				.rstn(rstn),
				.a0(P0450),
				.a1(P0460),
				.a2(P0470),
				.a3(P0550),
				.a4(P0560),
				.a5(P0570),
				.a6(P0650),
				.a7(P0660),
				.a8(P0670),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00451)
);

ninexnine_unit ninexnine_unit_772(
				.clk(clk),
				.rstn(rstn),
				.a0(P0451),
				.a1(P0461),
				.a2(P0471),
				.a3(P0551),
				.a4(P0561),
				.a5(P0571),
				.a6(P0651),
				.a7(P0661),
				.a8(P0671),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01451)
);

ninexnine_unit ninexnine_unit_773(
				.clk(clk),
				.rstn(rstn),
				.a0(P0452),
				.a1(P0462),
				.a2(P0472),
				.a3(P0552),
				.a4(P0562),
				.a5(P0572),
				.a6(P0652),
				.a7(P0662),
				.a8(P0672),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02451)
);

assign C0451=c00451+c01451+c02451;
assign A0451=(C0451>=0)?1:0;

ninexnine_unit ninexnine_unit_774(
				.clk(clk),
				.rstn(rstn),
				.a0(P0460),
				.a1(P0470),
				.a2(P0480),
				.a3(P0560),
				.a4(P0570),
				.a5(P0580),
				.a6(P0660),
				.a7(P0670),
				.a8(P0680),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00461)
);

ninexnine_unit ninexnine_unit_775(
				.clk(clk),
				.rstn(rstn),
				.a0(P0461),
				.a1(P0471),
				.a2(P0481),
				.a3(P0561),
				.a4(P0571),
				.a5(P0581),
				.a6(P0661),
				.a7(P0671),
				.a8(P0681),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01461)
);

ninexnine_unit ninexnine_unit_776(
				.clk(clk),
				.rstn(rstn),
				.a0(P0462),
				.a1(P0472),
				.a2(P0482),
				.a3(P0562),
				.a4(P0572),
				.a5(P0582),
				.a6(P0662),
				.a7(P0672),
				.a8(P0682),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02461)
);

assign C0461=c00461+c01461+c02461;
assign A0461=(C0461>=0)?1:0;

ninexnine_unit ninexnine_unit_777(
				.clk(clk),
				.rstn(rstn),
				.a0(P0470),
				.a1(P0480),
				.a2(P0490),
				.a3(P0570),
				.a4(P0580),
				.a5(P0590),
				.a6(P0670),
				.a7(P0680),
				.a8(P0690),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00471)
);

ninexnine_unit ninexnine_unit_778(
				.clk(clk),
				.rstn(rstn),
				.a0(P0471),
				.a1(P0481),
				.a2(P0491),
				.a3(P0571),
				.a4(P0581),
				.a5(P0591),
				.a6(P0671),
				.a7(P0681),
				.a8(P0691),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01471)
);

ninexnine_unit ninexnine_unit_779(
				.clk(clk),
				.rstn(rstn),
				.a0(P0472),
				.a1(P0482),
				.a2(P0492),
				.a3(P0572),
				.a4(P0582),
				.a5(P0592),
				.a6(P0672),
				.a7(P0682),
				.a8(P0692),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02471)
);

assign C0471=c00471+c01471+c02471;
assign A0471=(C0471>=0)?1:0;

ninexnine_unit ninexnine_unit_780(
				.clk(clk),
				.rstn(rstn),
				.a0(P0480),
				.a1(P0490),
				.a2(P04A0),
				.a3(P0580),
				.a4(P0590),
				.a5(P05A0),
				.a6(P0680),
				.a7(P0690),
				.a8(P06A0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00481)
);

ninexnine_unit ninexnine_unit_781(
				.clk(clk),
				.rstn(rstn),
				.a0(P0481),
				.a1(P0491),
				.a2(P04A1),
				.a3(P0581),
				.a4(P0591),
				.a5(P05A1),
				.a6(P0681),
				.a7(P0691),
				.a8(P06A1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01481)
);

ninexnine_unit ninexnine_unit_782(
				.clk(clk),
				.rstn(rstn),
				.a0(P0482),
				.a1(P0492),
				.a2(P04A2),
				.a3(P0582),
				.a4(P0592),
				.a5(P05A2),
				.a6(P0682),
				.a7(P0692),
				.a8(P06A2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02481)
);

assign C0481=c00481+c01481+c02481;
assign A0481=(C0481>=0)?1:0;

ninexnine_unit ninexnine_unit_783(
				.clk(clk),
				.rstn(rstn),
				.a0(P0490),
				.a1(P04A0),
				.a2(P04B0),
				.a3(P0590),
				.a4(P05A0),
				.a5(P05B0),
				.a6(P0690),
				.a7(P06A0),
				.a8(P06B0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00491)
);

ninexnine_unit ninexnine_unit_784(
				.clk(clk),
				.rstn(rstn),
				.a0(P0491),
				.a1(P04A1),
				.a2(P04B1),
				.a3(P0591),
				.a4(P05A1),
				.a5(P05B1),
				.a6(P0691),
				.a7(P06A1),
				.a8(P06B1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01491)
);

ninexnine_unit ninexnine_unit_785(
				.clk(clk),
				.rstn(rstn),
				.a0(P0492),
				.a1(P04A2),
				.a2(P04B2),
				.a3(P0592),
				.a4(P05A2),
				.a5(P05B2),
				.a6(P0692),
				.a7(P06A2),
				.a8(P06B2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02491)
);

assign C0491=c00491+c01491+c02491;
assign A0491=(C0491>=0)?1:0;

ninexnine_unit ninexnine_unit_786(
				.clk(clk),
				.rstn(rstn),
				.a0(P04A0),
				.a1(P04B0),
				.a2(P04C0),
				.a3(P05A0),
				.a4(P05B0),
				.a5(P05C0),
				.a6(P06A0),
				.a7(P06B0),
				.a8(P06C0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c004A1)
);

ninexnine_unit ninexnine_unit_787(
				.clk(clk),
				.rstn(rstn),
				.a0(P04A1),
				.a1(P04B1),
				.a2(P04C1),
				.a3(P05A1),
				.a4(P05B1),
				.a5(P05C1),
				.a6(P06A1),
				.a7(P06B1),
				.a8(P06C1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c014A1)
);

ninexnine_unit ninexnine_unit_788(
				.clk(clk),
				.rstn(rstn),
				.a0(P04A2),
				.a1(P04B2),
				.a2(P04C2),
				.a3(P05A2),
				.a4(P05B2),
				.a5(P05C2),
				.a6(P06A2),
				.a7(P06B2),
				.a8(P06C2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c024A1)
);

assign C04A1=c004A1+c014A1+c024A1;
assign A04A1=(C04A1>=0)?1:0;

ninexnine_unit ninexnine_unit_789(
				.clk(clk),
				.rstn(rstn),
				.a0(P04B0),
				.a1(P04C0),
				.a2(P04D0),
				.a3(P05B0),
				.a4(P05C0),
				.a5(P05D0),
				.a6(P06B0),
				.a7(P06C0),
				.a8(P06D0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c004B1)
);

ninexnine_unit ninexnine_unit_790(
				.clk(clk),
				.rstn(rstn),
				.a0(P04B1),
				.a1(P04C1),
				.a2(P04D1),
				.a3(P05B1),
				.a4(P05C1),
				.a5(P05D1),
				.a6(P06B1),
				.a7(P06C1),
				.a8(P06D1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c014B1)
);

ninexnine_unit ninexnine_unit_791(
				.clk(clk),
				.rstn(rstn),
				.a0(P04B2),
				.a1(P04C2),
				.a2(P04D2),
				.a3(P05B2),
				.a4(P05C2),
				.a5(P05D2),
				.a6(P06B2),
				.a7(P06C2),
				.a8(P06D2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c024B1)
);

assign C04B1=c004B1+c014B1+c024B1;
assign A04B1=(C04B1>=0)?1:0;

ninexnine_unit ninexnine_unit_792(
				.clk(clk),
				.rstn(rstn),
				.a0(P04C0),
				.a1(P04D0),
				.a2(P04E0),
				.a3(P05C0),
				.a4(P05D0),
				.a5(P05E0),
				.a6(P06C0),
				.a7(P06D0),
				.a8(P06E0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c004C1)
);

ninexnine_unit ninexnine_unit_793(
				.clk(clk),
				.rstn(rstn),
				.a0(P04C1),
				.a1(P04D1),
				.a2(P04E1),
				.a3(P05C1),
				.a4(P05D1),
				.a5(P05E1),
				.a6(P06C1),
				.a7(P06D1),
				.a8(P06E1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c014C1)
);

ninexnine_unit ninexnine_unit_794(
				.clk(clk),
				.rstn(rstn),
				.a0(P04C2),
				.a1(P04D2),
				.a2(P04E2),
				.a3(P05C2),
				.a4(P05D2),
				.a5(P05E2),
				.a6(P06C2),
				.a7(P06D2),
				.a8(P06E2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c024C1)
);

assign C04C1=c004C1+c014C1+c024C1;
assign A04C1=(C04C1>=0)?1:0;

ninexnine_unit ninexnine_unit_795(
				.clk(clk),
				.rstn(rstn),
				.a0(P04D0),
				.a1(P04E0),
				.a2(P04F0),
				.a3(P05D0),
				.a4(P05E0),
				.a5(P05F0),
				.a6(P06D0),
				.a7(P06E0),
				.a8(P06F0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c004D1)
);

ninexnine_unit ninexnine_unit_796(
				.clk(clk),
				.rstn(rstn),
				.a0(P04D1),
				.a1(P04E1),
				.a2(P04F1),
				.a3(P05D1),
				.a4(P05E1),
				.a5(P05F1),
				.a6(P06D1),
				.a7(P06E1),
				.a8(P06F1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c014D1)
);

ninexnine_unit ninexnine_unit_797(
				.clk(clk),
				.rstn(rstn),
				.a0(P04D2),
				.a1(P04E2),
				.a2(P04F2),
				.a3(P05D2),
				.a4(P05E2),
				.a5(P05F2),
				.a6(P06D2),
				.a7(P06E2),
				.a8(P06F2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c024D1)
);

assign C04D1=c004D1+c014D1+c024D1;
assign A04D1=(C04D1>=0)?1:0;

ninexnine_unit ninexnine_unit_798(
				.clk(clk),
				.rstn(rstn),
				.a0(P0500),
				.a1(P0510),
				.a2(P0520),
				.a3(P0600),
				.a4(P0610),
				.a5(P0620),
				.a6(P0700),
				.a7(P0710),
				.a8(P0720),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00501)
);

ninexnine_unit ninexnine_unit_799(
				.clk(clk),
				.rstn(rstn),
				.a0(P0501),
				.a1(P0511),
				.a2(P0521),
				.a3(P0601),
				.a4(P0611),
				.a5(P0621),
				.a6(P0701),
				.a7(P0711),
				.a8(P0721),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01501)
);

ninexnine_unit ninexnine_unit_800(
				.clk(clk),
				.rstn(rstn),
				.a0(P0502),
				.a1(P0512),
				.a2(P0522),
				.a3(P0602),
				.a4(P0612),
				.a5(P0622),
				.a6(P0702),
				.a7(P0712),
				.a8(P0722),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02501)
);

assign C0501=c00501+c01501+c02501;
assign A0501=(C0501>=0)?1:0;

ninexnine_unit ninexnine_unit_801(
				.clk(clk),
				.rstn(rstn),
				.a0(P0510),
				.a1(P0520),
				.a2(P0530),
				.a3(P0610),
				.a4(P0620),
				.a5(P0630),
				.a6(P0710),
				.a7(P0720),
				.a8(P0730),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00511)
);

ninexnine_unit ninexnine_unit_802(
				.clk(clk),
				.rstn(rstn),
				.a0(P0511),
				.a1(P0521),
				.a2(P0531),
				.a3(P0611),
				.a4(P0621),
				.a5(P0631),
				.a6(P0711),
				.a7(P0721),
				.a8(P0731),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01511)
);

ninexnine_unit ninexnine_unit_803(
				.clk(clk),
				.rstn(rstn),
				.a0(P0512),
				.a1(P0522),
				.a2(P0532),
				.a3(P0612),
				.a4(P0622),
				.a5(P0632),
				.a6(P0712),
				.a7(P0722),
				.a8(P0732),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02511)
);

assign C0511=c00511+c01511+c02511;
assign A0511=(C0511>=0)?1:0;

ninexnine_unit ninexnine_unit_804(
				.clk(clk),
				.rstn(rstn),
				.a0(P0520),
				.a1(P0530),
				.a2(P0540),
				.a3(P0620),
				.a4(P0630),
				.a5(P0640),
				.a6(P0720),
				.a7(P0730),
				.a8(P0740),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00521)
);

ninexnine_unit ninexnine_unit_805(
				.clk(clk),
				.rstn(rstn),
				.a0(P0521),
				.a1(P0531),
				.a2(P0541),
				.a3(P0621),
				.a4(P0631),
				.a5(P0641),
				.a6(P0721),
				.a7(P0731),
				.a8(P0741),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01521)
);

ninexnine_unit ninexnine_unit_806(
				.clk(clk),
				.rstn(rstn),
				.a0(P0522),
				.a1(P0532),
				.a2(P0542),
				.a3(P0622),
				.a4(P0632),
				.a5(P0642),
				.a6(P0722),
				.a7(P0732),
				.a8(P0742),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02521)
);

assign C0521=c00521+c01521+c02521;
assign A0521=(C0521>=0)?1:0;

ninexnine_unit ninexnine_unit_807(
				.clk(clk),
				.rstn(rstn),
				.a0(P0530),
				.a1(P0540),
				.a2(P0550),
				.a3(P0630),
				.a4(P0640),
				.a5(P0650),
				.a6(P0730),
				.a7(P0740),
				.a8(P0750),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00531)
);

ninexnine_unit ninexnine_unit_808(
				.clk(clk),
				.rstn(rstn),
				.a0(P0531),
				.a1(P0541),
				.a2(P0551),
				.a3(P0631),
				.a4(P0641),
				.a5(P0651),
				.a6(P0731),
				.a7(P0741),
				.a8(P0751),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01531)
);

ninexnine_unit ninexnine_unit_809(
				.clk(clk),
				.rstn(rstn),
				.a0(P0532),
				.a1(P0542),
				.a2(P0552),
				.a3(P0632),
				.a4(P0642),
				.a5(P0652),
				.a6(P0732),
				.a7(P0742),
				.a8(P0752),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02531)
);

assign C0531=c00531+c01531+c02531;
assign A0531=(C0531>=0)?1:0;

ninexnine_unit ninexnine_unit_810(
				.clk(clk),
				.rstn(rstn),
				.a0(P0540),
				.a1(P0550),
				.a2(P0560),
				.a3(P0640),
				.a4(P0650),
				.a5(P0660),
				.a6(P0740),
				.a7(P0750),
				.a8(P0760),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00541)
);

ninexnine_unit ninexnine_unit_811(
				.clk(clk),
				.rstn(rstn),
				.a0(P0541),
				.a1(P0551),
				.a2(P0561),
				.a3(P0641),
				.a4(P0651),
				.a5(P0661),
				.a6(P0741),
				.a7(P0751),
				.a8(P0761),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01541)
);

ninexnine_unit ninexnine_unit_812(
				.clk(clk),
				.rstn(rstn),
				.a0(P0542),
				.a1(P0552),
				.a2(P0562),
				.a3(P0642),
				.a4(P0652),
				.a5(P0662),
				.a6(P0742),
				.a7(P0752),
				.a8(P0762),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02541)
);

assign C0541=c00541+c01541+c02541;
assign A0541=(C0541>=0)?1:0;

ninexnine_unit ninexnine_unit_813(
				.clk(clk),
				.rstn(rstn),
				.a0(P0550),
				.a1(P0560),
				.a2(P0570),
				.a3(P0650),
				.a4(P0660),
				.a5(P0670),
				.a6(P0750),
				.a7(P0760),
				.a8(P0770),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00551)
);

ninexnine_unit ninexnine_unit_814(
				.clk(clk),
				.rstn(rstn),
				.a0(P0551),
				.a1(P0561),
				.a2(P0571),
				.a3(P0651),
				.a4(P0661),
				.a5(P0671),
				.a6(P0751),
				.a7(P0761),
				.a8(P0771),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01551)
);

ninexnine_unit ninexnine_unit_815(
				.clk(clk),
				.rstn(rstn),
				.a0(P0552),
				.a1(P0562),
				.a2(P0572),
				.a3(P0652),
				.a4(P0662),
				.a5(P0672),
				.a6(P0752),
				.a7(P0762),
				.a8(P0772),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02551)
);

assign C0551=c00551+c01551+c02551;
assign A0551=(C0551>=0)?1:0;

ninexnine_unit ninexnine_unit_816(
				.clk(clk),
				.rstn(rstn),
				.a0(P0560),
				.a1(P0570),
				.a2(P0580),
				.a3(P0660),
				.a4(P0670),
				.a5(P0680),
				.a6(P0760),
				.a7(P0770),
				.a8(P0780),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00561)
);

ninexnine_unit ninexnine_unit_817(
				.clk(clk),
				.rstn(rstn),
				.a0(P0561),
				.a1(P0571),
				.a2(P0581),
				.a3(P0661),
				.a4(P0671),
				.a5(P0681),
				.a6(P0761),
				.a7(P0771),
				.a8(P0781),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01561)
);

ninexnine_unit ninexnine_unit_818(
				.clk(clk),
				.rstn(rstn),
				.a0(P0562),
				.a1(P0572),
				.a2(P0582),
				.a3(P0662),
				.a4(P0672),
				.a5(P0682),
				.a6(P0762),
				.a7(P0772),
				.a8(P0782),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02561)
);

assign C0561=c00561+c01561+c02561;
assign A0561=(C0561>=0)?1:0;

ninexnine_unit ninexnine_unit_819(
				.clk(clk),
				.rstn(rstn),
				.a0(P0570),
				.a1(P0580),
				.a2(P0590),
				.a3(P0670),
				.a4(P0680),
				.a5(P0690),
				.a6(P0770),
				.a7(P0780),
				.a8(P0790),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00571)
);

ninexnine_unit ninexnine_unit_820(
				.clk(clk),
				.rstn(rstn),
				.a0(P0571),
				.a1(P0581),
				.a2(P0591),
				.a3(P0671),
				.a4(P0681),
				.a5(P0691),
				.a6(P0771),
				.a7(P0781),
				.a8(P0791),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01571)
);

ninexnine_unit ninexnine_unit_821(
				.clk(clk),
				.rstn(rstn),
				.a0(P0572),
				.a1(P0582),
				.a2(P0592),
				.a3(P0672),
				.a4(P0682),
				.a5(P0692),
				.a6(P0772),
				.a7(P0782),
				.a8(P0792),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02571)
);

assign C0571=c00571+c01571+c02571;
assign A0571=(C0571>=0)?1:0;

ninexnine_unit ninexnine_unit_822(
				.clk(clk),
				.rstn(rstn),
				.a0(P0580),
				.a1(P0590),
				.a2(P05A0),
				.a3(P0680),
				.a4(P0690),
				.a5(P06A0),
				.a6(P0780),
				.a7(P0790),
				.a8(P07A0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00581)
);

ninexnine_unit ninexnine_unit_823(
				.clk(clk),
				.rstn(rstn),
				.a0(P0581),
				.a1(P0591),
				.a2(P05A1),
				.a3(P0681),
				.a4(P0691),
				.a5(P06A1),
				.a6(P0781),
				.a7(P0791),
				.a8(P07A1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01581)
);

ninexnine_unit ninexnine_unit_824(
				.clk(clk),
				.rstn(rstn),
				.a0(P0582),
				.a1(P0592),
				.a2(P05A2),
				.a3(P0682),
				.a4(P0692),
				.a5(P06A2),
				.a6(P0782),
				.a7(P0792),
				.a8(P07A2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02581)
);

assign C0581=c00581+c01581+c02581;
assign A0581=(C0581>=0)?1:0;

ninexnine_unit ninexnine_unit_825(
				.clk(clk),
				.rstn(rstn),
				.a0(P0590),
				.a1(P05A0),
				.a2(P05B0),
				.a3(P0690),
				.a4(P06A0),
				.a5(P06B0),
				.a6(P0790),
				.a7(P07A0),
				.a8(P07B0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00591)
);

ninexnine_unit ninexnine_unit_826(
				.clk(clk),
				.rstn(rstn),
				.a0(P0591),
				.a1(P05A1),
				.a2(P05B1),
				.a3(P0691),
				.a4(P06A1),
				.a5(P06B1),
				.a6(P0791),
				.a7(P07A1),
				.a8(P07B1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01591)
);

ninexnine_unit ninexnine_unit_827(
				.clk(clk),
				.rstn(rstn),
				.a0(P0592),
				.a1(P05A2),
				.a2(P05B2),
				.a3(P0692),
				.a4(P06A2),
				.a5(P06B2),
				.a6(P0792),
				.a7(P07A2),
				.a8(P07B2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02591)
);

assign C0591=c00591+c01591+c02591;
assign A0591=(C0591>=0)?1:0;

ninexnine_unit ninexnine_unit_828(
				.clk(clk),
				.rstn(rstn),
				.a0(P05A0),
				.a1(P05B0),
				.a2(P05C0),
				.a3(P06A0),
				.a4(P06B0),
				.a5(P06C0),
				.a6(P07A0),
				.a7(P07B0),
				.a8(P07C0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c005A1)
);

ninexnine_unit ninexnine_unit_829(
				.clk(clk),
				.rstn(rstn),
				.a0(P05A1),
				.a1(P05B1),
				.a2(P05C1),
				.a3(P06A1),
				.a4(P06B1),
				.a5(P06C1),
				.a6(P07A1),
				.a7(P07B1),
				.a8(P07C1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c015A1)
);

ninexnine_unit ninexnine_unit_830(
				.clk(clk),
				.rstn(rstn),
				.a0(P05A2),
				.a1(P05B2),
				.a2(P05C2),
				.a3(P06A2),
				.a4(P06B2),
				.a5(P06C2),
				.a6(P07A2),
				.a7(P07B2),
				.a8(P07C2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c025A1)
);

assign C05A1=c005A1+c015A1+c025A1;
assign A05A1=(C05A1>=0)?1:0;

ninexnine_unit ninexnine_unit_831(
				.clk(clk),
				.rstn(rstn),
				.a0(P05B0),
				.a1(P05C0),
				.a2(P05D0),
				.a3(P06B0),
				.a4(P06C0),
				.a5(P06D0),
				.a6(P07B0),
				.a7(P07C0),
				.a8(P07D0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c005B1)
);

ninexnine_unit ninexnine_unit_832(
				.clk(clk),
				.rstn(rstn),
				.a0(P05B1),
				.a1(P05C1),
				.a2(P05D1),
				.a3(P06B1),
				.a4(P06C1),
				.a5(P06D1),
				.a6(P07B1),
				.a7(P07C1),
				.a8(P07D1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c015B1)
);

ninexnine_unit ninexnine_unit_833(
				.clk(clk),
				.rstn(rstn),
				.a0(P05B2),
				.a1(P05C2),
				.a2(P05D2),
				.a3(P06B2),
				.a4(P06C2),
				.a5(P06D2),
				.a6(P07B2),
				.a7(P07C2),
				.a8(P07D2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c025B1)
);

assign C05B1=c005B1+c015B1+c025B1;
assign A05B1=(C05B1>=0)?1:0;

ninexnine_unit ninexnine_unit_834(
				.clk(clk),
				.rstn(rstn),
				.a0(P05C0),
				.a1(P05D0),
				.a2(P05E0),
				.a3(P06C0),
				.a4(P06D0),
				.a5(P06E0),
				.a6(P07C0),
				.a7(P07D0),
				.a8(P07E0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c005C1)
);

ninexnine_unit ninexnine_unit_835(
				.clk(clk),
				.rstn(rstn),
				.a0(P05C1),
				.a1(P05D1),
				.a2(P05E1),
				.a3(P06C1),
				.a4(P06D1),
				.a5(P06E1),
				.a6(P07C1),
				.a7(P07D1),
				.a8(P07E1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c015C1)
);

ninexnine_unit ninexnine_unit_836(
				.clk(clk),
				.rstn(rstn),
				.a0(P05C2),
				.a1(P05D2),
				.a2(P05E2),
				.a3(P06C2),
				.a4(P06D2),
				.a5(P06E2),
				.a6(P07C2),
				.a7(P07D2),
				.a8(P07E2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c025C1)
);

assign C05C1=c005C1+c015C1+c025C1;
assign A05C1=(C05C1>=0)?1:0;

ninexnine_unit ninexnine_unit_837(
				.clk(clk),
				.rstn(rstn),
				.a0(P05D0),
				.a1(P05E0),
				.a2(P05F0),
				.a3(P06D0),
				.a4(P06E0),
				.a5(P06F0),
				.a6(P07D0),
				.a7(P07E0),
				.a8(P07F0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c005D1)
);

ninexnine_unit ninexnine_unit_838(
				.clk(clk),
				.rstn(rstn),
				.a0(P05D1),
				.a1(P05E1),
				.a2(P05F1),
				.a3(P06D1),
				.a4(P06E1),
				.a5(P06F1),
				.a6(P07D1),
				.a7(P07E1),
				.a8(P07F1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c015D1)
);

ninexnine_unit ninexnine_unit_839(
				.clk(clk),
				.rstn(rstn),
				.a0(P05D2),
				.a1(P05E2),
				.a2(P05F2),
				.a3(P06D2),
				.a4(P06E2),
				.a5(P06F2),
				.a6(P07D2),
				.a7(P07E2),
				.a8(P07F2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c025D1)
);

assign C05D1=c005D1+c015D1+c025D1;
assign A05D1=(C05D1>=0)?1:0;

ninexnine_unit ninexnine_unit_840(
				.clk(clk),
				.rstn(rstn),
				.a0(P0600),
				.a1(P0610),
				.a2(P0620),
				.a3(P0700),
				.a4(P0710),
				.a5(P0720),
				.a6(P0800),
				.a7(P0810),
				.a8(P0820),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00601)
);

ninexnine_unit ninexnine_unit_841(
				.clk(clk),
				.rstn(rstn),
				.a0(P0601),
				.a1(P0611),
				.a2(P0621),
				.a3(P0701),
				.a4(P0711),
				.a5(P0721),
				.a6(P0801),
				.a7(P0811),
				.a8(P0821),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01601)
);

ninexnine_unit ninexnine_unit_842(
				.clk(clk),
				.rstn(rstn),
				.a0(P0602),
				.a1(P0612),
				.a2(P0622),
				.a3(P0702),
				.a4(P0712),
				.a5(P0722),
				.a6(P0802),
				.a7(P0812),
				.a8(P0822),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02601)
);

assign C0601=c00601+c01601+c02601;
assign A0601=(C0601>=0)?1:0;

ninexnine_unit ninexnine_unit_843(
				.clk(clk),
				.rstn(rstn),
				.a0(P0610),
				.a1(P0620),
				.a2(P0630),
				.a3(P0710),
				.a4(P0720),
				.a5(P0730),
				.a6(P0810),
				.a7(P0820),
				.a8(P0830),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00611)
);

ninexnine_unit ninexnine_unit_844(
				.clk(clk),
				.rstn(rstn),
				.a0(P0611),
				.a1(P0621),
				.a2(P0631),
				.a3(P0711),
				.a4(P0721),
				.a5(P0731),
				.a6(P0811),
				.a7(P0821),
				.a8(P0831),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01611)
);

ninexnine_unit ninexnine_unit_845(
				.clk(clk),
				.rstn(rstn),
				.a0(P0612),
				.a1(P0622),
				.a2(P0632),
				.a3(P0712),
				.a4(P0722),
				.a5(P0732),
				.a6(P0812),
				.a7(P0822),
				.a8(P0832),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02611)
);

assign C0611=c00611+c01611+c02611;
assign A0611=(C0611>=0)?1:0;

ninexnine_unit ninexnine_unit_846(
				.clk(clk),
				.rstn(rstn),
				.a0(P0620),
				.a1(P0630),
				.a2(P0640),
				.a3(P0720),
				.a4(P0730),
				.a5(P0740),
				.a6(P0820),
				.a7(P0830),
				.a8(P0840),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00621)
);

ninexnine_unit ninexnine_unit_847(
				.clk(clk),
				.rstn(rstn),
				.a0(P0621),
				.a1(P0631),
				.a2(P0641),
				.a3(P0721),
				.a4(P0731),
				.a5(P0741),
				.a6(P0821),
				.a7(P0831),
				.a8(P0841),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01621)
);

ninexnine_unit ninexnine_unit_848(
				.clk(clk),
				.rstn(rstn),
				.a0(P0622),
				.a1(P0632),
				.a2(P0642),
				.a3(P0722),
				.a4(P0732),
				.a5(P0742),
				.a6(P0822),
				.a7(P0832),
				.a8(P0842),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02621)
);

assign C0621=c00621+c01621+c02621;
assign A0621=(C0621>=0)?1:0;

ninexnine_unit ninexnine_unit_849(
				.clk(clk),
				.rstn(rstn),
				.a0(P0630),
				.a1(P0640),
				.a2(P0650),
				.a3(P0730),
				.a4(P0740),
				.a5(P0750),
				.a6(P0830),
				.a7(P0840),
				.a8(P0850),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00631)
);

ninexnine_unit ninexnine_unit_850(
				.clk(clk),
				.rstn(rstn),
				.a0(P0631),
				.a1(P0641),
				.a2(P0651),
				.a3(P0731),
				.a4(P0741),
				.a5(P0751),
				.a6(P0831),
				.a7(P0841),
				.a8(P0851),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01631)
);

ninexnine_unit ninexnine_unit_851(
				.clk(clk),
				.rstn(rstn),
				.a0(P0632),
				.a1(P0642),
				.a2(P0652),
				.a3(P0732),
				.a4(P0742),
				.a5(P0752),
				.a6(P0832),
				.a7(P0842),
				.a8(P0852),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02631)
);

assign C0631=c00631+c01631+c02631;
assign A0631=(C0631>=0)?1:0;

ninexnine_unit ninexnine_unit_852(
				.clk(clk),
				.rstn(rstn),
				.a0(P0640),
				.a1(P0650),
				.a2(P0660),
				.a3(P0740),
				.a4(P0750),
				.a5(P0760),
				.a6(P0840),
				.a7(P0850),
				.a8(P0860),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00641)
);

ninexnine_unit ninexnine_unit_853(
				.clk(clk),
				.rstn(rstn),
				.a0(P0641),
				.a1(P0651),
				.a2(P0661),
				.a3(P0741),
				.a4(P0751),
				.a5(P0761),
				.a6(P0841),
				.a7(P0851),
				.a8(P0861),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01641)
);

ninexnine_unit ninexnine_unit_854(
				.clk(clk),
				.rstn(rstn),
				.a0(P0642),
				.a1(P0652),
				.a2(P0662),
				.a3(P0742),
				.a4(P0752),
				.a5(P0762),
				.a6(P0842),
				.a7(P0852),
				.a8(P0862),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02641)
);

assign C0641=c00641+c01641+c02641;
assign A0641=(C0641>=0)?1:0;

ninexnine_unit ninexnine_unit_855(
				.clk(clk),
				.rstn(rstn),
				.a0(P0650),
				.a1(P0660),
				.a2(P0670),
				.a3(P0750),
				.a4(P0760),
				.a5(P0770),
				.a6(P0850),
				.a7(P0860),
				.a8(P0870),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00651)
);

ninexnine_unit ninexnine_unit_856(
				.clk(clk),
				.rstn(rstn),
				.a0(P0651),
				.a1(P0661),
				.a2(P0671),
				.a3(P0751),
				.a4(P0761),
				.a5(P0771),
				.a6(P0851),
				.a7(P0861),
				.a8(P0871),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01651)
);

ninexnine_unit ninexnine_unit_857(
				.clk(clk),
				.rstn(rstn),
				.a0(P0652),
				.a1(P0662),
				.a2(P0672),
				.a3(P0752),
				.a4(P0762),
				.a5(P0772),
				.a6(P0852),
				.a7(P0862),
				.a8(P0872),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02651)
);

assign C0651=c00651+c01651+c02651;
assign A0651=(C0651>=0)?1:0;

ninexnine_unit ninexnine_unit_858(
				.clk(clk),
				.rstn(rstn),
				.a0(P0660),
				.a1(P0670),
				.a2(P0680),
				.a3(P0760),
				.a4(P0770),
				.a5(P0780),
				.a6(P0860),
				.a7(P0870),
				.a8(P0880),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00661)
);

ninexnine_unit ninexnine_unit_859(
				.clk(clk),
				.rstn(rstn),
				.a0(P0661),
				.a1(P0671),
				.a2(P0681),
				.a3(P0761),
				.a4(P0771),
				.a5(P0781),
				.a6(P0861),
				.a7(P0871),
				.a8(P0881),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01661)
);

ninexnine_unit ninexnine_unit_860(
				.clk(clk),
				.rstn(rstn),
				.a0(P0662),
				.a1(P0672),
				.a2(P0682),
				.a3(P0762),
				.a4(P0772),
				.a5(P0782),
				.a6(P0862),
				.a7(P0872),
				.a8(P0882),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02661)
);

assign C0661=c00661+c01661+c02661;
assign A0661=(C0661>=0)?1:0;

ninexnine_unit ninexnine_unit_861(
				.clk(clk),
				.rstn(rstn),
				.a0(P0670),
				.a1(P0680),
				.a2(P0690),
				.a3(P0770),
				.a4(P0780),
				.a5(P0790),
				.a6(P0870),
				.a7(P0880),
				.a8(P0890),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00671)
);

ninexnine_unit ninexnine_unit_862(
				.clk(clk),
				.rstn(rstn),
				.a0(P0671),
				.a1(P0681),
				.a2(P0691),
				.a3(P0771),
				.a4(P0781),
				.a5(P0791),
				.a6(P0871),
				.a7(P0881),
				.a8(P0891),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01671)
);

ninexnine_unit ninexnine_unit_863(
				.clk(clk),
				.rstn(rstn),
				.a0(P0672),
				.a1(P0682),
				.a2(P0692),
				.a3(P0772),
				.a4(P0782),
				.a5(P0792),
				.a6(P0872),
				.a7(P0882),
				.a8(P0892),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02671)
);

assign C0671=c00671+c01671+c02671;
assign A0671=(C0671>=0)?1:0;

ninexnine_unit ninexnine_unit_864(
				.clk(clk),
				.rstn(rstn),
				.a0(P0680),
				.a1(P0690),
				.a2(P06A0),
				.a3(P0780),
				.a4(P0790),
				.a5(P07A0),
				.a6(P0880),
				.a7(P0890),
				.a8(P08A0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00681)
);

ninexnine_unit ninexnine_unit_865(
				.clk(clk),
				.rstn(rstn),
				.a0(P0681),
				.a1(P0691),
				.a2(P06A1),
				.a3(P0781),
				.a4(P0791),
				.a5(P07A1),
				.a6(P0881),
				.a7(P0891),
				.a8(P08A1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01681)
);

ninexnine_unit ninexnine_unit_866(
				.clk(clk),
				.rstn(rstn),
				.a0(P0682),
				.a1(P0692),
				.a2(P06A2),
				.a3(P0782),
				.a4(P0792),
				.a5(P07A2),
				.a6(P0882),
				.a7(P0892),
				.a8(P08A2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02681)
);

assign C0681=c00681+c01681+c02681;
assign A0681=(C0681>=0)?1:0;

ninexnine_unit ninexnine_unit_867(
				.clk(clk),
				.rstn(rstn),
				.a0(P0690),
				.a1(P06A0),
				.a2(P06B0),
				.a3(P0790),
				.a4(P07A0),
				.a5(P07B0),
				.a6(P0890),
				.a7(P08A0),
				.a8(P08B0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00691)
);

ninexnine_unit ninexnine_unit_868(
				.clk(clk),
				.rstn(rstn),
				.a0(P0691),
				.a1(P06A1),
				.a2(P06B1),
				.a3(P0791),
				.a4(P07A1),
				.a5(P07B1),
				.a6(P0891),
				.a7(P08A1),
				.a8(P08B1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01691)
);

ninexnine_unit ninexnine_unit_869(
				.clk(clk),
				.rstn(rstn),
				.a0(P0692),
				.a1(P06A2),
				.a2(P06B2),
				.a3(P0792),
				.a4(P07A2),
				.a5(P07B2),
				.a6(P0892),
				.a7(P08A2),
				.a8(P08B2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02691)
);

assign C0691=c00691+c01691+c02691;
assign A0691=(C0691>=0)?1:0;

ninexnine_unit ninexnine_unit_870(
				.clk(clk),
				.rstn(rstn),
				.a0(P06A0),
				.a1(P06B0),
				.a2(P06C0),
				.a3(P07A0),
				.a4(P07B0),
				.a5(P07C0),
				.a6(P08A0),
				.a7(P08B0),
				.a8(P08C0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c006A1)
);

ninexnine_unit ninexnine_unit_871(
				.clk(clk),
				.rstn(rstn),
				.a0(P06A1),
				.a1(P06B1),
				.a2(P06C1),
				.a3(P07A1),
				.a4(P07B1),
				.a5(P07C1),
				.a6(P08A1),
				.a7(P08B1),
				.a8(P08C1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c016A1)
);

ninexnine_unit ninexnine_unit_872(
				.clk(clk),
				.rstn(rstn),
				.a0(P06A2),
				.a1(P06B2),
				.a2(P06C2),
				.a3(P07A2),
				.a4(P07B2),
				.a5(P07C2),
				.a6(P08A2),
				.a7(P08B2),
				.a8(P08C2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c026A1)
);

assign C06A1=c006A1+c016A1+c026A1;
assign A06A1=(C06A1>=0)?1:0;

ninexnine_unit ninexnine_unit_873(
				.clk(clk),
				.rstn(rstn),
				.a0(P06B0),
				.a1(P06C0),
				.a2(P06D0),
				.a3(P07B0),
				.a4(P07C0),
				.a5(P07D0),
				.a6(P08B0),
				.a7(P08C0),
				.a8(P08D0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c006B1)
);

ninexnine_unit ninexnine_unit_874(
				.clk(clk),
				.rstn(rstn),
				.a0(P06B1),
				.a1(P06C1),
				.a2(P06D1),
				.a3(P07B1),
				.a4(P07C1),
				.a5(P07D1),
				.a6(P08B1),
				.a7(P08C1),
				.a8(P08D1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c016B1)
);

ninexnine_unit ninexnine_unit_875(
				.clk(clk),
				.rstn(rstn),
				.a0(P06B2),
				.a1(P06C2),
				.a2(P06D2),
				.a3(P07B2),
				.a4(P07C2),
				.a5(P07D2),
				.a6(P08B2),
				.a7(P08C2),
				.a8(P08D2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c026B1)
);

assign C06B1=c006B1+c016B1+c026B1;
assign A06B1=(C06B1>=0)?1:0;

ninexnine_unit ninexnine_unit_876(
				.clk(clk),
				.rstn(rstn),
				.a0(P06C0),
				.a1(P06D0),
				.a2(P06E0),
				.a3(P07C0),
				.a4(P07D0),
				.a5(P07E0),
				.a6(P08C0),
				.a7(P08D0),
				.a8(P08E0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c006C1)
);

ninexnine_unit ninexnine_unit_877(
				.clk(clk),
				.rstn(rstn),
				.a0(P06C1),
				.a1(P06D1),
				.a2(P06E1),
				.a3(P07C1),
				.a4(P07D1),
				.a5(P07E1),
				.a6(P08C1),
				.a7(P08D1),
				.a8(P08E1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c016C1)
);

ninexnine_unit ninexnine_unit_878(
				.clk(clk),
				.rstn(rstn),
				.a0(P06C2),
				.a1(P06D2),
				.a2(P06E2),
				.a3(P07C2),
				.a4(P07D2),
				.a5(P07E2),
				.a6(P08C2),
				.a7(P08D2),
				.a8(P08E2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c026C1)
);

assign C06C1=c006C1+c016C1+c026C1;
assign A06C1=(C06C1>=0)?1:0;

ninexnine_unit ninexnine_unit_879(
				.clk(clk),
				.rstn(rstn),
				.a0(P06D0),
				.a1(P06E0),
				.a2(P06F0),
				.a3(P07D0),
				.a4(P07E0),
				.a5(P07F0),
				.a6(P08D0),
				.a7(P08E0),
				.a8(P08F0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c006D1)
);

ninexnine_unit ninexnine_unit_880(
				.clk(clk),
				.rstn(rstn),
				.a0(P06D1),
				.a1(P06E1),
				.a2(P06F1),
				.a3(P07D1),
				.a4(P07E1),
				.a5(P07F1),
				.a6(P08D1),
				.a7(P08E1),
				.a8(P08F1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c016D1)
);

ninexnine_unit ninexnine_unit_881(
				.clk(clk),
				.rstn(rstn),
				.a0(P06D2),
				.a1(P06E2),
				.a2(P06F2),
				.a3(P07D2),
				.a4(P07E2),
				.a5(P07F2),
				.a6(P08D2),
				.a7(P08E2),
				.a8(P08F2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c026D1)
);

assign C06D1=c006D1+c016D1+c026D1;
assign A06D1=(C06D1>=0)?1:0;

ninexnine_unit ninexnine_unit_882(
				.clk(clk),
				.rstn(rstn),
				.a0(P0700),
				.a1(P0710),
				.a2(P0720),
				.a3(P0800),
				.a4(P0810),
				.a5(P0820),
				.a6(P0900),
				.a7(P0910),
				.a8(P0920),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00701)
);

ninexnine_unit ninexnine_unit_883(
				.clk(clk),
				.rstn(rstn),
				.a0(P0701),
				.a1(P0711),
				.a2(P0721),
				.a3(P0801),
				.a4(P0811),
				.a5(P0821),
				.a6(P0901),
				.a7(P0911),
				.a8(P0921),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01701)
);

ninexnine_unit ninexnine_unit_884(
				.clk(clk),
				.rstn(rstn),
				.a0(P0702),
				.a1(P0712),
				.a2(P0722),
				.a3(P0802),
				.a4(P0812),
				.a5(P0822),
				.a6(P0902),
				.a7(P0912),
				.a8(P0922),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02701)
);

assign C0701=c00701+c01701+c02701;
assign A0701=(C0701>=0)?1:0;

ninexnine_unit ninexnine_unit_885(
				.clk(clk),
				.rstn(rstn),
				.a0(P0710),
				.a1(P0720),
				.a2(P0730),
				.a3(P0810),
				.a4(P0820),
				.a5(P0830),
				.a6(P0910),
				.a7(P0920),
				.a8(P0930),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00711)
);

ninexnine_unit ninexnine_unit_886(
				.clk(clk),
				.rstn(rstn),
				.a0(P0711),
				.a1(P0721),
				.a2(P0731),
				.a3(P0811),
				.a4(P0821),
				.a5(P0831),
				.a6(P0911),
				.a7(P0921),
				.a8(P0931),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01711)
);

ninexnine_unit ninexnine_unit_887(
				.clk(clk),
				.rstn(rstn),
				.a0(P0712),
				.a1(P0722),
				.a2(P0732),
				.a3(P0812),
				.a4(P0822),
				.a5(P0832),
				.a6(P0912),
				.a7(P0922),
				.a8(P0932),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02711)
);

assign C0711=c00711+c01711+c02711;
assign A0711=(C0711>=0)?1:0;

ninexnine_unit ninexnine_unit_888(
				.clk(clk),
				.rstn(rstn),
				.a0(P0720),
				.a1(P0730),
				.a2(P0740),
				.a3(P0820),
				.a4(P0830),
				.a5(P0840),
				.a6(P0920),
				.a7(P0930),
				.a8(P0940),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00721)
);

ninexnine_unit ninexnine_unit_889(
				.clk(clk),
				.rstn(rstn),
				.a0(P0721),
				.a1(P0731),
				.a2(P0741),
				.a3(P0821),
				.a4(P0831),
				.a5(P0841),
				.a6(P0921),
				.a7(P0931),
				.a8(P0941),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01721)
);

ninexnine_unit ninexnine_unit_890(
				.clk(clk),
				.rstn(rstn),
				.a0(P0722),
				.a1(P0732),
				.a2(P0742),
				.a3(P0822),
				.a4(P0832),
				.a5(P0842),
				.a6(P0922),
				.a7(P0932),
				.a8(P0942),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02721)
);

assign C0721=c00721+c01721+c02721;
assign A0721=(C0721>=0)?1:0;

ninexnine_unit ninexnine_unit_891(
				.clk(clk),
				.rstn(rstn),
				.a0(P0730),
				.a1(P0740),
				.a2(P0750),
				.a3(P0830),
				.a4(P0840),
				.a5(P0850),
				.a6(P0930),
				.a7(P0940),
				.a8(P0950),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00731)
);

ninexnine_unit ninexnine_unit_892(
				.clk(clk),
				.rstn(rstn),
				.a0(P0731),
				.a1(P0741),
				.a2(P0751),
				.a3(P0831),
				.a4(P0841),
				.a5(P0851),
				.a6(P0931),
				.a7(P0941),
				.a8(P0951),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01731)
);

ninexnine_unit ninexnine_unit_893(
				.clk(clk),
				.rstn(rstn),
				.a0(P0732),
				.a1(P0742),
				.a2(P0752),
				.a3(P0832),
				.a4(P0842),
				.a5(P0852),
				.a6(P0932),
				.a7(P0942),
				.a8(P0952),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02731)
);

assign C0731=c00731+c01731+c02731;
assign A0731=(C0731>=0)?1:0;

ninexnine_unit ninexnine_unit_894(
				.clk(clk),
				.rstn(rstn),
				.a0(P0740),
				.a1(P0750),
				.a2(P0760),
				.a3(P0840),
				.a4(P0850),
				.a5(P0860),
				.a6(P0940),
				.a7(P0950),
				.a8(P0960),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00741)
);

ninexnine_unit ninexnine_unit_895(
				.clk(clk),
				.rstn(rstn),
				.a0(P0741),
				.a1(P0751),
				.a2(P0761),
				.a3(P0841),
				.a4(P0851),
				.a5(P0861),
				.a6(P0941),
				.a7(P0951),
				.a8(P0961),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01741)
);

ninexnine_unit ninexnine_unit_896(
				.clk(clk),
				.rstn(rstn),
				.a0(P0742),
				.a1(P0752),
				.a2(P0762),
				.a3(P0842),
				.a4(P0852),
				.a5(P0862),
				.a6(P0942),
				.a7(P0952),
				.a8(P0962),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02741)
);

assign C0741=c00741+c01741+c02741;
assign A0741=(C0741>=0)?1:0;

ninexnine_unit ninexnine_unit_897(
				.clk(clk),
				.rstn(rstn),
				.a0(P0750),
				.a1(P0760),
				.a2(P0770),
				.a3(P0850),
				.a4(P0860),
				.a5(P0870),
				.a6(P0950),
				.a7(P0960),
				.a8(P0970),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00751)
);

ninexnine_unit ninexnine_unit_898(
				.clk(clk),
				.rstn(rstn),
				.a0(P0751),
				.a1(P0761),
				.a2(P0771),
				.a3(P0851),
				.a4(P0861),
				.a5(P0871),
				.a6(P0951),
				.a7(P0961),
				.a8(P0971),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01751)
);

ninexnine_unit ninexnine_unit_899(
				.clk(clk),
				.rstn(rstn),
				.a0(P0752),
				.a1(P0762),
				.a2(P0772),
				.a3(P0852),
				.a4(P0862),
				.a5(P0872),
				.a6(P0952),
				.a7(P0962),
				.a8(P0972),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02751)
);

assign C0751=c00751+c01751+c02751;
assign A0751=(C0751>=0)?1:0;

ninexnine_unit ninexnine_unit_900(
				.clk(clk),
				.rstn(rstn),
				.a0(P0760),
				.a1(P0770),
				.a2(P0780),
				.a3(P0860),
				.a4(P0870),
				.a5(P0880),
				.a6(P0960),
				.a7(P0970),
				.a8(P0980),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00761)
);

ninexnine_unit ninexnine_unit_901(
				.clk(clk),
				.rstn(rstn),
				.a0(P0761),
				.a1(P0771),
				.a2(P0781),
				.a3(P0861),
				.a4(P0871),
				.a5(P0881),
				.a6(P0961),
				.a7(P0971),
				.a8(P0981),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01761)
);

ninexnine_unit ninexnine_unit_902(
				.clk(clk),
				.rstn(rstn),
				.a0(P0762),
				.a1(P0772),
				.a2(P0782),
				.a3(P0862),
				.a4(P0872),
				.a5(P0882),
				.a6(P0962),
				.a7(P0972),
				.a8(P0982),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02761)
);

assign C0761=c00761+c01761+c02761;
assign A0761=(C0761>=0)?1:0;

ninexnine_unit ninexnine_unit_903(
				.clk(clk),
				.rstn(rstn),
				.a0(P0770),
				.a1(P0780),
				.a2(P0790),
				.a3(P0870),
				.a4(P0880),
				.a5(P0890),
				.a6(P0970),
				.a7(P0980),
				.a8(P0990),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00771)
);

ninexnine_unit ninexnine_unit_904(
				.clk(clk),
				.rstn(rstn),
				.a0(P0771),
				.a1(P0781),
				.a2(P0791),
				.a3(P0871),
				.a4(P0881),
				.a5(P0891),
				.a6(P0971),
				.a7(P0981),
				.a8(P0991),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01771)
);

ninexnine_unit ninexnine_unit_905(
				.clk(clk),
				.rstn(rstn),
				.a0(P0772),
				.a1(P0782),
				.a2(P0792),
				.a3(P0872),
				.a4(P0882),
				.a5(P0892),
				.a6(P0972),
				.a7(P0982),
				.a8(P0992),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02771)
);

assign C0771=c00771+c01771+c02771;
assign A0771=(C0771>=0)?1:0;

ninexnine_unit ninexnine_unit_906(
				.clk(clk),
				.rstn(rstn),
				.a0(P0780),
				.a1(P0790),
				.a2(P07A0),
				.a3(P0880),
				.a4(P0890),
				.a5(P08A0),
				.a6(P0980),
				.a7(P0990),
				.a8(P09A0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00781)
);

ninexnine_unit ninexnine_unit_907(
				.clk(clk),
				.rstn(rstn),
				.a0(P0781),
				.a1(P0791),
				.a2(P07A1),
				.a3(P0881),
				.a4(P0891),
				.a5(P08A1),
				.a6(P0981),
				.a7(P0991),
				.a8(P09A1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01781)
);

ninexnine_unit ninexnine_unit_908(
				.clk(clk),
				.rstn(rstn),
				.a0(P0782),
				.a1(P0792),
				.a2(P07A2),
				.a3(P0882),
				.a4(P0892),
				.a5(P08A2),
				.a6(P0982),
				.a7(P0992),
				.a8(P09A2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02781)
);

assign C0781=c00781+c01781+c02781;
assign A0781=(C0781>=0)?1:0;

ninexnine_unit ninexnine_unit_909(
				.clk(clk),
				.rstn(rstn),
				.a0(P0790),
				.a1(P07A0),
				.a2(P07B0),
				.a3(P0890),
				.a4(P08A0),
				.a5(P08B0),
				.a6(P0990),
				.a7(P09A0),
				.a8(P09B0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00791)
);

ninexnine_unit ninexnine_unit_910(
				.clk(clk),
				.rstn(rstn),
				.a0(P0791),
				.a1(P07A1),
				.a2(P07B1),
				.a3(P0891),
				.a4(P08A1),
				.a5(P08B1),
				.a6(P0991),
				.a7(P09A1),
				.a8(P09B1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01791)
);

ninexnine_unit ninexnine_unit_911(
				.clk(clk),
				.rstn(rstn),
				.a0(P0792),
				.a1(P07A2),
				.a2(P07B2),
				.a3(P0892),
				.a4(P08A2),
				.a5(P08B2),
				.a6(P0992),
				.a7(P09A2),
				.a8(P09B2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02791)
);

assign C0791=c00791+c01791+c02791;
assign A0791=(C0791>=0)?1:0;

ninexnine_unit ninexnine_unit_912(
				.clk(clk),
				.rstn(rstn),
				.a0(P07A0),
				.a1(P07B0),
				.a2(P07C0),
				.a3(P08A0),
				.a4(P08B0),
				.a5(P08C0),
				.a6(P09A0),
				.a7(P09B0),
				.a8(P09C0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c007A1)
);

ninexnine_unit ninexnine_unit_913(
				.clk(clk),
				.rstn(rstn),
				.a0(P07A1),
				.a1(P07B1),
				.a2(P07C1),
				.a3(P08A1),
				.a4(P08B1),
				.a5(P08C1),
				.a6(P09A1),
				.a7(P09B1),
				.a8(P09C1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c017A1)
);

ninexnine_unit ninexnine_unit_914(
				.clk(clk),
				.rstn(rstn),
				.a0(P07A2),
				.a1(P07B2),
				.a2(P07C2),
				.a3(P08A2),
				.a4(P08B2),
				.a5(P08C2),
				.a6(P09A2),
				.a7(P09B2),
				.a8(P09C2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c027A1)
);

assign C07A1=c007A1+c017A1+c027A1;
assign A07A1=(C07A1>=0)?1:0;

ninexnine_unit ninexnine_unit_915(
				.clk(clk),
				.rstn(rstn),
				.a0(P07B0),
				.a1(P07C0),
				.a2(P07D0),
				.a3(P08B0),
				.a4(P08C0),
				.a5(P08D0),
				.a6(P09B0),
				.a7(P09C0),
				.a8(P09D0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c007B1)
);

ninexnine_unit ninexnine_unit_916(
				.clk(clk),
				.rstn(rstn),
				.a0(P07B1),
				.a1(P07C1),
				.a2(P07D1),
				.a3(P08B1),
				.a4(P08C1),
				.a5(P08D1),
				.a6(P09B1),
				.a7(P09C1),
				.a8(P09D1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c017B1)
);

ninexnine_unit ninexnine_unit_917(
				.clk(clk),
				.rstn(rstn),
				.a0(P07B2),
				.a1(P07C2),
				.a2(P07D2),
				.a3(P08B2),
				.a4(P08C2),
				.a5(P08D2),
				.a6(P09B2),
				.a7(P09C2),
				.a8(P09D2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c027B1)
);

assign C07B1=c007B1+c017B1+c027B1;
assign A07B1=(C07B1>=0)?1:0;

ninexnine_unit ninexnine_unit_918(
				.clk(clk),
				.rstn(rstn),
				.a0(P07C0),
				.a1(P07D0),
				.a2(P07E0),
				.a3(P08C0),
				.a4(P08D0),
				.a5(P08E0),
				.a6(P09C0),
				.a7(P09D0),
				.a8(P09E0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c007C1)
);

ninexnine_unit ninexnine_unit_919(
				.clk(clk),
				.rstn(rstn),
				.a0(P07C1),
				.a1(P07D1),
				.a2(P07E1),
				.a3(P08C1),
				.a4(P08D1),
				.a5(P08E1),
				.a6(P09C1),
				.a7(P09D1),
				.a8(P09E1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c017C1)
);

ninexnine_unit ninexnine_unit_920(
				.clk(clk),
				.rstn(rstn),
				.a0(P07C2),
				.a1(P07D2),
				.a2(P07E2),
				.a3(P08C2),
				.a4(P08D2),
				.a5(P08E2),
				.a6(P09C2),
				.a7(P09D2),
				.a8(P09E2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c027C1)
);

assign C07C1=c007C1+c017C1+c027C1;
assign A07C1=(C07C1>=0)?1:0;

ninexnine_unit ninexnine_unit_921(
				.clk(clk),
				.rstn(rstn),
				.a0(P07D0),
				.a1(P07E0),
				.a2(P07F0),
				.a3(P08D0),
				.a4(P08E0),
				.a5(P08F0),
				.a6(P09D0),
				.a7(P09E0),
				.a8(P09F0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c007D1)
);

ninexnine_unit ninexnine_unit_922(
				.clk(clk),
				.rstn(rstn),
				.a0(P07D1),
				.a1(P07E1),
				.a2(P07F1),
				.a3(P08D1),
				.a4(P08E1),
				.a5(P08F1),
				.a6(P09D1),
				.a7(P09E1),
				.a8(P09F1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c017D1)
);

ninexnine_unit ninexnine_unit_923(
				.clk(clk),
				.rstn(rstn),
				.a0(P07D2),
				.a1(P07E2),
				.a2(P07F2),
				.a3(P08D2),
				.a4(P08E2),
				.a5(P08F2),
				.a6(P09D2),
				.a7(P09E2),
				.a8(P09F2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c027D1)
);

assign C07D1=c007D1+c017D1+c027D1;
assign A07D1=(C07D1>=0)?1:0;

ninexnine_unit ninexnine_unit_924(
				.clk(clk),
				.rstn(rstn),
				.a0(P0800),
				.a1(P0810),
				.a2(P0820),
				.a3(P0900),
				.a4(P0910),
				.a5(P0920),
				.a6(P0A00),
				.a7(P0A10),
				.a8(P0A20),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00801)
);

ninexnine_unit ninexnine_unit_925(
				.clk(clk),
				.rstn(rstn),
				.a0(P0801),
				.a1(P0811),
				.a2(P0821),
				.a3(P0901),
				.a4(P0911),
				.a5(P0921),
				.a6(P0A01),
				.a7(P0A11),
				.a8(P0A21),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01801)
);

ninexnine_unit ninexnine_unit_926(
				.clk(clk),
				.rstn(rstn),
				.a0(P0802),
				.a1(P0812),
				.a2(P0822),
				.a3(P0902),
				.a4(P0912),
				.a5(P0922),
				.a6(P0A02),
				.a7(P0A12),
				.a8(P0A22),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02801)
);

assign C0801=c00801+c01801+c02801;
assign A0801=(C0801>=0)?1:0;

ninexnine_unit ninexnine_unit_927(
				.clk(clk),
				.rstn(rstn),
				.a0(P0810),
				.a1(P0820),
				.a2(P0830),
				.a3(P0910),
				.a4(P0920),
				.a5(P0930),
				.a6(P0A10),
				.a7(P0A20),
				.a8(P0A30),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00811)
);

ninexnine_unit ninexnine_unit_928(
				.clk(clk),
				.rstn(rstn),
				.a0(P0811),
				.a1(P0821),
				.a2(P0831),
				.a3(P0911),
				.a4(P0921),
				.a5(P0931),
				.a6(P0A11),
				.a7(P0A21),
				.a8(P0A31),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01811)
);

ninexnine_unit ninexnine_unit_929(
				.clk(clk),
				.rstn(rstn),
				.a0(P0812),
				.a1(P0822),
				.a2(P0832),
				.a3(P0912),
				.a4(P0922),
				.a5(P0932),
				.a6(P0A12),
				.a7(P0A22),
				.a8(P0A32),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02811)
);

assign C0811=c00811+c01811+c02811;
assign A0811=(C0811>=0)?1:0;

ninexnine_unit ninexnine_unit_930(
				.clk(clk),
				.rstn(rstn),
				.a0(P0820),
				.a1(P0830),
				.a2(P0840),
				.a3(P0920),
				.a4(P0930),
				.a5(P0940),
				.a6(P0A20),
				.a7(P0A30),
				.a8(P0A40),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00821)
);

ninexnine_unit ninexnine_unit_931(
				.clk(clk),
				.rstn(rstn),
				.a0(P0821),
				.a1(P0831),
				.a2(P0841),
				.a3(P0921),
				.a4(P0931),
				.a5(P0941),
				.a6(P0A21),
				.a7(P0A31),
				.a8(P0A41),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01821)
);

ninexnine_unit ninexnine_unit_932(
				.clk(clk),
				.rstn(rstn),
				.a0(P0822),
				.a1(P0832),
				.a2(P0842),
				.a3(P0922),
				.a4(P0932),
				.a5(P0942),
				.a6(P0A22),
				.a7(P0A32),
				.a8(P0A42),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02821)
);

assign C0821=c00821+c01821+c02821;
assign A0821=(C0821>=0)?1:0;

ninexnine_unit ninexnine_unit_933(
				.clk(clk),
				.rstn(rstn),
				.a0(P0830),
				.a1(P0840),
				.a2(P0850),
				.a3(P0930),
				.a4(P0940),
				.a5(P0950),
				.a6(P0A30),
				.a7(P0A40),
				.a8(P0A50),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00831)
);

ninexnine_unit ninexnine_unit_934(
				.clk(clk),
				.rstn(rstn),
				.a0(P0831),
				.a1(P0841),
				.a2(P0851),
				.a3(P0931),
				.a4(P0941),
				.a5(P0951),
				.a6(P0A31),
				.a7(P0A41),
				.a8(P0A51),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01831)
);

ninexnine_unit ninexnine_unit_935(
				.clk(clk),
				.rstn(rstn),
				.a0(P0832),
				.a1(P0842),
				.a2(P0852),
				.a3(P0932),
				.a4(P0942),
				.a5(P0952),
				.a6(P0A32),
				.a7(P0A42),
				.a8(P0A52),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02831)
);

assign C0831=c00831+c01831+c02831;
assign A0831=(C0831>=0)?1:0;

ninexnine_unit ninexnine_unit_936(
				.clk(clk),
				.rstn(rstn),
				.a0(P0840),
				.a1(P0850),
				.a2(P0860),
				.a3(P0940),
				.a4(P0950),
				.a5(P0960),
				.a6(P0A40),
				.a7(P0A50),
				.a8(P0A60),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00841)
);

ninexnine_unit ninexnine_unit_937(
				.clk(clk),
				.rstn(rstn),
				.a0(P0841),
				.a1(P0851),
				.a2(P0861),
				.a3(P0941),
				.a4(P0951),
				.a5(P0961),
				.a6(P0A41),
				.a7(P0A51),
				.a8(P0A61),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01841)
);

ninexnine_unit ninexnine_unit_938(
				.clk(clk),
				.rstn(rstn),
				.a0(P0842),
				.a1(P0852),
				.a2(P0862),
				.a3(P0942),
				.a4(P0952),
				.a5(P0962),
				.a6(P0A42),
				.a7(P0A52),
				.a8(P0A62),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02841)
);

assign C0841=c00841+c01841+c02841;
assign A0841=(C0841>=0)?1:0;

ninexnine_unit ninexnine_unit_939(
				.clk(clk),
				.rstn(rstn),
				.a0(P0850),
				.a1(P0860),
				.a2(P0870),
				.a3(P0950),
				.a4(P0960),
				.a5(P0970),
				.a6(P0A50),
				.a7(P0A60),
				.a8(P0A70),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00851)
);

ninexnine_unit ninexnine_unit_940(
				.clk(clk),
				.rstn(rstn),
				.a0(P0851),
				.a1(P0861),
				.a2(P0871),
				.a3(P0951),
				.a4(P0961),
				.a5(P0971),
				.a6(P0A51),
				.a7(P0A61),
				.a8(P0A71),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01851)
);

ninexnine_unit ninexnine_unit_941(
				.clk(clk),
				.rstn(rstn),
				.a0(P0852),
				.a1(P0862),
				.a2(P0872),
				.a3(P0952),
				.a4(P0962),
				.a5(P0972),
				.a6(P0A52),
				.a7(P0A62),
				.a8(P0A72),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02851)
);

assign C0851=c00851+c01851+c02851;
assign A0851=(C0851>=0)?1:0;

ninexnine_unit ninexnine_unit_942(
				.clk(clk),
				.rstn(rstn),
				.a0(P0860),
				.a1(P0870),
				.a2(P0880),
				.a3(P0960),
				.a4(P0970),
				.a5(P0980),
				.a6(P0A60),
				.a7(P0A70),
				.a8(P0A80),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00861)
);

ninexnine_unit ninexnine_unit_943(
				.clk(clk),
				.rstn(rstn),
				.a0(P0861),
				.a1(P0871),
				.a2(P0881),
				.a3(P0961),
				.a4(P0971),
				.a5(P0981),
				.a6(P0A61),
				.a7(P0A71),
				.a8(P0A81),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01861)
);

ninexnine_unit ninexnine_unit_944(
				.clk(clk),
				.rstn(rstn),
				.a0(P0862),
				.a1(P0872),
				.a2(P0882),
				.a3(P0962),
				.a4(P0972),
				.a5(P0982),
				.a6(P0A62),
				.a7(P0A72),
				.a8(P0A82),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02861)
);

assign C0861=c00861+c01861+c02861;
assign A0861=(C0861>=0)?1:0;

ninexnine_unit ninexnine_unit_945(
				.clk(clk),
				.rstn(rstn),
				.a0(P0870),
				.a1(P0880),
				.a2(P0890),
				.a3(P0970),
				.a4(P0980),
				.a5(P0990),
				.a6(P0A70),
				.a7(P0A80),
				.a8(P0A90),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00871)
);

ninexnine_unit ninexnine_unit_946(
				.clk(clk),
				.rstn(rstn),
				.a0(P0871),
				.a1(P0881),
				.a2(P0891),
				.a3(P0971),
				.a4(P0981),
				.a5(P0991),
				.a6(P0A71),
				.a7(P0A81),
				.a8(P0A91),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01871)
);

ninexnine_unit ninexnine_unit_947(
				.clk(clk),
				.rstn(rstn),
				.a0(P0872),
				.a1(P0882),
				.a2(P0892),
				.a3(P0972),
				.a4(P0982),
				.a5(P0992),
				.a6(P0A72),
				.a7(P0A82),
				.a8(P0A92),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02871)
);

assign C0871=c00871+c01871+c02871;
assign A0871=(C0871>=0)?1:0;

ninexnine_unit ninexnine_unit_948(
				.clk(clk),
				.rstn(rstn),
				.a0(P0880),
				.a1(P0890),
				.a2(P08A0),
				.a3(P0980),
				.a4(P0990),
				.a5(P09A0),
				.a6(P0A80),
				.a7(P0A90),
				.a8(P0AA0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00881)
);

ninexnine_unit ninexnine_unit_949(
				.clk(clk),
				.rstn(rstn),
				.a0(P0881),
				.a1(P0891),
				.a2(P08A1),
				.a3(P0981),
				.a4(P0991),
				.a5(P09A1),
				.a6(P0A81),
				.a7(P0A91),
				.a8(P0AA1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01881)
);

ninexnine_unit ninexnine_unit_950(
				.clk(clk),
				.rstn(rstn),
				.a0(P0882),
				.a1(P0892),
				.a2(P08A2),
				.a3(P0982),
				.a4(P0992),
				.a5(P09A2),
				.a6(P0A82),
				.a7(P0A92),
				.a8(P0AA2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02881)
);

assign C0881=c00881+c01881+c02881;
assign A0881=(C0881>=0)?1:0;

ninexnine_unit ninexnine_unit_951(
				.clk(clk),
				.rstn(rstn),
				.a0(P0890),
				.a1(P08A0),
				.a2(P08B0),
				.a3(P0990),
				.a4(P09A0),
				.a5(P09B0),
				.a6(P0A90),
				.a7(P0AA0),
				.a8(P0AB0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00891)
);

ninexnine_unit ninexnine_unit_952(
				.clk(clk),
				.rstn(rstn),
				.a0(P0891),
				.a1(P08A1),
				.a2(P08B1),
				.a3(P0991),
				.a4(P09A1),
				.a5(P09B1),
				.a6(P0A91),
				.a7(P0AA1),
				.a8(P0AB1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01891)
);

ninexnine_unit ninexnine_unit_953(
				.clk(clk),
				.rstn(rstn),
				.a0(P0892),
				.a1(P08A2),
				.a2(P08B2),
				.a3(P0992),
				.a4(P09A2),
				.a5(P09B2),
				.a6(P0A92),
				.a7(P0AA2),
				.a8(P0AB2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02891)
);

assign C0891=c00891+c01891+c02891;
assign A0891=(C0891>=0)?1:0;

ninexnine_unit ninexnine_unit_954(
				.clk(clk),
				.rstn(rstn),
				.a0(P08A0),
				.a1(P08B0),
				.a2(P08C0),
				.a3(P09A0),
				.a4(P09B0),
				.a5(P09C0),
				.a6(P0AA0),
				.a7(P0AB0),
				.a8(P0AC0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c008A1)
);

ninexnine_unit ninexnine_unit_955(
				.clk(clk),
				.rstn(rstn),
				.a0(P08A1),
				.a1(P08B1),
				.a2(P08C1),
				.a3(P09A1),
				.a4(P09B1),
				.a5(P09C1),
				.a6(P0AA1),
				.a7(P0AB1),
				.a8(P0AC1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c018A1)
);

ninexnine_unit ninexnine_unit_956(
				.clk(clk),
				.rstn(rstn),
				.a0(P08A2),
				.a1(P08B2),
				.a2(P08C2),
				.a3(P09A2),
				.a4(P09B2),
				.a5(P09C2),
				.a6(P0AA2),
				.a7(P0AB2),
				.a8(P0AC2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c028A1)
);

assign C08A1=c008A1+c018A1+c028A1;
assign A08A1=(C08A1>=0)?1:0;

ninexnine_unit ninexnine_unit_957(
				.clk(clk),
				.rstn(rstn),
				.a0(P08B0),
				.a1(P08C0),
				.a2(P08D0),
				.a3(P09B0),
				.a4(P09C0),
				.a5(P09D0),
				.a6(P0AB0),
				.a7(P0AC0),
				.a8(P0AD0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c008B1)
);

ninexnine_unit ninexnine_unit_958(
				.clk(clk),
				.rstn(rstn),
				.a0(P08B1),
				.a1(P08C1),
				.a2(P08D1),
				.a3(P09B1),
				.a4(P09C1),
				.a5(P09D1),
				.a6(P0AB1),
				.a7(P0AC1),
				.a8(P0AD1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c018B1)
);

ninexnine_unit ninexnine_unit_959(
				.clk(clk),
				.rstn(rstn),
				.a0(P08B2),
				.a1(P08C2),
				.a2(P08D2),
				.a3(P09B2),
				.a4(P09C2),
				.a5(P09D2),
				.a6(P0AB2),
				.a7(P0AC2),
				.a8(P0AD2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c028B1)
);

assign C08B1=c008B1+c018B1+c028B1;
assign A08B1=(C08B1>=0)?1:0;

ninexnine_unit ninexnine_unit_960(
				.clk(clk),
				.rstn(rstn),
				.a0(P08C0),
				.a1(P08D0),
				.a2(P08E0),
				.a3(P09C0),
				.a4(P09D0),
				.a5(P09E0),
				.a6(P0AC0),
				.a7(P0AD0),
				.a8(P0AE0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c008C1)
);

ninexnine_unit ninexnine_unit_961(
				.clk(clk),
				.rstn(rstn),
				.a0(P08C1),
				.a1(P08D1),
				.a2(P08E1),
				.a3(P09C1),
				.a4(P09D1),
				.a5(P09E1),
				.a6(P0AC1),
				.a7(P0AD1),
				.a8(P0AE1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c018C1)
);

ninexnine_unit ninexnine_unit_962(
				.clk(clk),
				.rstn(rstn),
				.a0(P08C2),
				.a1(P08D2),
				.a2(P08E2),
				.a3(P09C2),
				.a4(P09D2),
				.a5(P09E2),
				.a6(P0AC2),
				.a7(P0AD2),
				.a8(P0AE2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c028C1)
);

assign C08C1=c008C1+c018C1+c028C1;
assign A08C1=(C08C1>=0)?1:0;

ninexnine_unit ninexnine_unit_963(
				.clk(clk),
				.rstn(rstn),
				.a0(P08D0),
				.a1(P08E0),
				.a2(P08F0),
				.a3(P09D0),
				.a4(P09E0),
				.a5(P09F0),
				.a6(P0AD0),
				.a7(P0AE0),
				.a8(P0AF0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c008D1)
);

ninexnine_unit ninexnine_unit_964(
				.clk(clk),
				.rstn(rstn),
				.a0(P08D1),
				.a1(P08E1),
				.a2(P08F1),
				.a3(P09D1),
				.a4(P09E1),
				.a5(P09F1),
				.a6(P0AD1),
				.a7(P0AE1),
				.a8(P0AF1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c018D1)
);

ninexnine_unit ninexnine_unit_965(
				.clk(clk),
				.rstn(rstn),
				.a0(P08D2),
				.a1(P08E2),
				.a2(P08F2),
				.a3(P09D2),
				.a4(P09E2),
				.a5(P09F2),
				.a6(P0AD2),
				.a7(P0AE2),
				.a8(P0AF2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c028D1)
);

assign C08D1=c008D1+c018D1+c028D1;
assign A08D1=(C08D1>=0)?1:0;

ninexnine_unit ninexnine_unit_966(
				.clk(clk),
				.rstn(rstn),
				.a0(P0900),
				.a1(P0910),
				.a2(P0920),
				.a3(P0A00),
				.a4(P0A10),
				.a5(P0A20),
				.a6(P0B00),
				.a7(P0B10),
				.a8(P0B20),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00901)
);

ninexnine_unit ninexnine_unit_967(
				.clk(clk),
				.rstn(rstn),
				.a0(P0901),
				.a1(P0911),
				.a2(P0921),
				.a3(P0A01),
				.a4(P0A11),
				.a5(P0A21),
				.a6(P0B01),
				.a7(P0B11),
				.a8(P0B21),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01901)
);

ninexnine_unit ninexnine_unit_968(
				.clk(clk),
				.rstn(rstn),
				.a0(P0902),
				.a1(P0912),
				.a2(P0922),
				.a3(P0A02),
				.a4(P0A12),
				.a5(P0A22),
				.a6(P0B02),
				.a7(P0B12),
				.a8(P0B22),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02901)
);

assign C0901=c00901+c01901+c02901;
assign A0901=(C0901>=0)?1:0;

ninexnine_unit ninexnine_unit_969(
				.clk(clk),
				.rstn(rstn),
				.a0(P0910),
				.a1(P0920),
				.a2(P0930),
				.a3(P0A10),
				.a4(P0A20),
				.a5(P0A30),
				.a6(P0B10),
				.a7(P0B20),
				.a8(P0B30),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00911)
);

ninexnine_unit ninexnine_unit_970(
				.clk(clk),
				.rstn(rstn),
				.a0(P0911),
				.a1(P0921),
				.a2(P0931),
				.a3(P0A11),
				.a4(P0A21),
				.a5(P0A31),
				.a6(P0B11),
				.a7(P0B21),
				.a8(P0B31),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01911)
);

ninexnine_unit ninexnine_unit_971(
				.clk(clk),
				.rstn(rstn),
				.a0(P0912),
				.a1(P0922),
				.a2(P0932),
				.a3(P0A12),
				.a4(P0A22),
				.a5(P0A32),
				.a6(P0B12),
				.a7(P0B22),
				.a8(P0B32),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02911)
);

assign C0911=c00911+c01911+c02911;
assign A0911=(C0911>=0)?1:0;

ninexnine_unit ninexnine_unit_972(
				.clk(clk),
				.rstn(rstn),
				.a0(P0920),
				.a1(P0930),
				.a2(P0940),
				.a3(P0A20),
				.a4(P0A30),
				.a5(P0A40),
				.a6(P0B20),
				.a7(P0B30),
				.a8(P0B40),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00921)
);

ninexnine_unit ninexnine_unit_973(
				.clk(clk),
				.rstn(rstn),
				.a0(P0921),
				.a1(P0931),
				.a2(P0941),
				.a3(P0A21),
				.a4(P0A31),
				.a5(P0A41),
				.a6(P0B21),
				.a7(P0B31),
				.a8(P0B41),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01921)
);

ninexnine_unit ninexnine_unit_974(
				.clk(clk),
				.rstn(rstn),
				.a0(P0922),
				.a1(P0932),
				.a2(P0942),
				.a3(P0A22),
				.a4(P0A32),
				.a5(P0A42),
				.a6(P0B22),
				.a7(P0B32),
				.a8(P0B42),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02921)
);

assign C0921=c00921+c01921+c02921;
assign A0921=(C0921>=0)?1:0;

ninexnine_unit ninexnine_unit_975(
				.clk(clk),
				.rstn(rstn),
				.a0(P0930),
				.a1(P0940),
				.a2(P0950),
				.a3(P0A30),
				.a4(P0A40),
				.a5(P0A50),
				.a6(P0B30),
				.a7(P0B40),
				.a8(P0B50),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00931)
);

ninexnine_unit ninexnine_unit_976(
				.clk(clk),
				.rstn(rstn),
				.a0(P0931),
				.a1(P0941),
				.a2(P0951),
				.a3(P0A31),
				.a4(P0A41),
				.a5(P0A51),
				.a6(P0B31),
				.a7(P0B41),
				.a8(P0B51),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01931)
);

ninexnine_unit ninexnine_unit_977(
				.clk(clk),
				.rstn(rstn),
				.a0(P0932),
				.a1(P0942),
				.a2(P0952),
				.a3(P0A32),
				.a4(P0A42),
				.a5(P0A52),
				.a6(P0B32),
				.a7(P0B42),
				.a8(P0B52),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02931)
);

assign C0931=c00931+c01931+c02931;
assign A0931=(C0931>=0)?1:0;

ninexnine_unit ninexnine_unit_978(
				.clk(clk),
				.rstn(rstn),
				.a0(P0940),
				.a1(P0950),
				.a2(P0960),
				.a3(P0A40),
				.a4(P0A50),
				.a5(P0A60),
				.a6(P0B40),
				.a7(P0B50),
				.a8(P0B60),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00941)
);

ninexnine_unit ninexnine_unit_979(
				.clk(clk),
				.rstn(rstn),
				.a0(P0941),
				.a1(P0951),
				.a2(P0961),
				.a3(P0A41),
				.a4(P0A51),
				.a5(P0A61),
				.a6(P0B41),
				.a7(P0B51),
				.a8(P0B61),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01941)
);

ninexnine_unit ninexnine_unit_980(
				.clk(clk),
				.rstn(rstn),
				.a0(P0942),
				.a1(P0952),
				.a2(P0962),
				.a3(P0A42),
				.a4(P0A52),
				.a5(P0A62),
				.a6(P0B42),
				.a7(P0B52),
				.a8(P0B62),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02941)
);

assign C0941=c00941+c01941+c02941;
assign A0941=(C0941>=0)?1:0;

ninexnine_unit ninexnine_unit_981(
				.clk(clk),
				.rstn(rstn),
				.a0(P0950),
				.a1(P0960),
				.a2(P0970),
				.a3(P0A50),
				.a4(P0A60),
				.a5(P0A70),
				.a6(P0B50),
				.a7(P0B60),
				.a8(P0B70),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00951)
);

ninexnine_unit ninexnine_unit_982(
				.clk(clk),
				.rstn(rstn),
				.a0(P0951),
				.a1(P0961),
				.a2(P0971),
				.a3(P0A51),
				.a4(P0A61),
				.a5(P0A71),
				.a6(P0B51),
				.a7(P0B61),
				.a8(P0B71),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01951)
);

ninexnine_unit ninexnine_unit_983(
				.clk(clk),
				.rstn(rstn),
				.a0(P0952),
				.a1(P0962),
				.a2(P0972),
				.a3(P0A52),
				.a4(P0A62),
				.a5(P0A72),
				.a6(P0B52),
				.a7(P0B62),
				.a8(P0B72),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02951)
);

assign C0951=c00951+c01951+c02951;
assign A0951=(C0951>=0)?1:0;

ninexnine_unit ninexnine_unit_984(
				.clk(clk),
				.rstn(rstn),
				.a0(P0960),
				.a1(P0970),
				.a2(P0980),
				.a3(P0A60),
				.a4(P0A70),
				.a5(P0A80),
				.a6(P0B60),
				.a7(P0B70),
				.a8(P0B80),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00961)
);

ninexnine_unit ninexnine_unit_985(
				.clk(clk),
				.rstn(rstn),
				.a0(P0961),
				.a1(P0971),
				.a2(P0981),
				.a3(P0A61),
				.a4(P0A71),
				.a5(P0A81),
				.a6(P0B61),
				.a7(P0B71),
				.a8(P0B81),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01961)
);

ninexnine_unit ninexnine_unit_986(
				.clk(clk),
				.rstn(rstn),
				.a0(P0962),
				.a1(P0972),
				.a2(P0982),
				.a3(P0A62),
				.a4(P0A72),
				.a5(P0A82),
				.a6(P0B62),
				.a7(P0B72),
				.a8(P0B82),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02961)
);

assign C0961=c00961+c01961+c02961;
assign A0961=(C0961>=0)?1:0;

ninexnine_unit ninexnine_unit_987(
				.clk(clk),
				.rstn(rstn),
				.a0(P0970),
				.a1(P0980),
				.a2(P0990),
				.a3(P0A70),
				.a4(P0A80),
				.a5(P0A90),
				.a6(P0B70),
				.a7(P0B80),
				.a8(P0B90),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00971)
);

ninexnine_unit ninexnine_unit_988(
				.clk(clk),
				.rstn(rstn),
				.a0(P0971),
				.a1(P0981),
				.a2(P0991),
				.a3(P0A71),
				.a4(P0A81),
				.a5(P0A91),
				.a6(P0B71),
				.a7(P0B81),
				.a8(P0B91),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01971)
);

ninexnine_unit ninexnine_unit_989(
				.clk(clk),
				.rstn(rstn),
				.a0(P0972),
				.a1(P0982),
				.a2(P0992),
				.a3(P0A72),
				.a4(P0A82),
				.a5(P0A92),
				.a6(P0B72),
				.a7(P0B82),
				.a8(P0B92),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02971)
);

assign C0971=c00971+c01971+c02971;
assign A0971=(C0971>=0)?1:0;

ninexnine_unit ninexnine_unit_990(
				.clk(clk),
				.rstn(rstn),
				.a0(P0980),
				.a1(P0990),
				.a2(P09A0),
				.a3(P0A80),
				.a4(P0A90),
				.a5(P0AA0),
				.a6(P0B80),
				.a7(P0B90),
				.a8(P0BA0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00981)
);

ninexnine_unit ninexnine_unit_991(
				.clk(clk),
				.rstn(rstn),
				.a0(P0981),
				.a1(P0991),
				.a2(P09A1),
				.a3(P0A81),
				.a4(P0A91),
				.a5(P0AA1),
				.a6(P0B81),
				.a7(P0B91),
				.a8(P0BA1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01981)
);

ninexnine_unit ninexnine_unit_992(
				.clk(clk),
				.rstn(rstn),
				.a0(P0982),
				.a1(P0992),
				.a2(P09A2),
				.a3(P0A82),
				.a4(P0A92),
				.a5(P0AA2),
				.a6(P0B82),
				.a7(P0B92),
				.a8(P0BA2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02981)
);

assign C0981=c00981+c01981+c02981;
assign A0981=(C0981>=0)?1:0;

ninexnine_unit ninexnine_unit_993(
				.clk(clk),
				.rstn(rstn),
				.a0(P0990),
				.a1(P09A0),
				.a2(P09B0),
				.a3(P0A90),
				.a4(P0AA0),
				.a5(P0AB0),
				.a6(P0B90),
				.a7(P0BA0),
				.a8(P0BB0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00991)
);

ninexnine_unit ninexnine_unit_994(
				.clk(clk),
				.rstn(rstn),
				.a0(P0991),
				.a1(P09A1),
				.a2(P09B1),
				.a3(P0A91),
				.a4(P0AA1),
				.a5(P0AB1),
				.a6(P0B91),
				.a7(P0BA1),
				.a8(P0BB1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01991)
);

ninexnine_unit ninexnine_unit_995(
				.clk(clk),
				.rstn(rstn),
				.a0(P0992),
				.a1(P09A2),
				.a2(P09B2),
				.a3(P0A92),
				.a4(P0AA2),
				.a5(P0AB2),
				.a6(P0B92),
				.a7(P0BA2),
				.a8(P0BB2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02991)
);

assign C0991=c00991+c01991+c02991;
assign A0991=(C0991>=0)?1:0;

ninexnine_unit ninexnine_unit_996(
				.clk(clk),
				.rstn(rstn),
				.a0(P09A0),
				.a1(P09B0),
				.a2(P09C0),
				.a3(P0AA0),
				.a4(P0AB0),
				.a5(P0AC0),
				.a6(P0BA0),
				.a7(P0BB0),
				.a8(P0BC0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c009A1)
);

ninexnine_unit ninexnine_unit_997(
				.clk(clk),
				.rstn(rstn),
				.a0(P09A1),
				.a1(P09B1),
				.a2(P09C1),
				.a3(P0AA1),
				.a4(P0AB1),
				.a5(P0AC1),
				.a6(P0BA1),
				.a7(P0BB1),
				.a8(P0BC1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c019A1)
);

ninexnine_unit ninexnine_unit_998(
				.clk(clk),
				.rstn(rstn),
				.a0(P09A2),
				.a1(P09B2),
				.a2(P09C2),
				.a3(P0AA2),
				.a4(P0AB2),
				.a5(P0AC2),
				.a6(P0BA2),
				.a7(P0BB2),
				.a8(P0BC2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c029A1)
);

assign C09A1=c009A1+c019A1+c029A1;
assign A09A1=(C09A1>=0)?1:0;

ninexnine_unit ninexnine_unit_999(
				.clk(clk),
				.rstn(rstn),
				.a0(P09B0),
				.a1(P09C0),
				.a2(P09D0),
				.a3(P0AB0),
				.a4(P0AC0),
				.a5(P0AD0),
				.a6(P0BB0),
				.a7(P0BC0),
				.a8(P0BD0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c009B1)
);

ninexnine_unit ninexnine_unit_1000(
				.clk(clk),
				.rstn(rstn),
				.a0(P09B1),
				.a1(P09C1),
				.a2(P09D1),
				.a3(P0AB1),
				.a4(P0AC1),
				.a5(P0AD1),
				.a6(P0BB1),
				.a7(P0BC1),
				.a8(P0BD1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c019B1)
);

ninexnine_unit ninexnine_unit_1001(
				.clk(clk),
				.rstn(rstn),
				.a0(P09B2),
				.a1(P09C2),
				.a2(P09D2),
				.a3(P0AB2),
				.a4(P0AC2),
				.a5(P0AD2),
				.a6(P0BB2),
				.a7(P0BC2),
				.a8(P0BD2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c029B1)
);

assign C09B1=c009B1+c019B1+c029B1;
assign A09B1=(C09B1>=0)?1:0;

ninexnine_unit ninexnine_unit_1002(
				.clk(clk),
				.rstn(rstn),
				.a0(P09C0),
				.a1(P09D0),
				.a2(P09E0),
				.a3(P0AC0),
				.a4(P0AD0),
				.a5(P0AE0),
				.a6(P0BC0),
				.a7(P0BD0),
				.a8(P0BE0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c009C1)
);

ninexnine_unit ninexnine_unit_1003(
				.clk(clk),
				.rstn(rstn),
				.a0(P09C1),
				.a1(P09D1),
				.a2(P09E1),
				.a3(P0AC1),
				.a4(P0AD1),
				.a5(P0AE1),
				.a6(P0BC1),
				.a7(P0BD1),
				.a8(P0BE1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c019C1)
);

ninexnine_unit ninexnine_unit_1004(
				.clk(clk),
				.rstn(rstn),
				.a0(P09C2),
				.a1(P09D2),
				.a2(P09E2),
				.a3(P0AC2),
				.a4(P0AD2),
				.a5(P0AE2),
				.a6(P0BC2),
				.a7(P0BD2),
				.a8(P0BE2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c029C1)
);

assign C09C1=c009C1+c019C1+c029C1;
assign A09C1=(C09C1>=0)?1:0;

ninexnine_unit ninexnine_unit_1005(
				.clk(clk),
				.rstn(rstn),
				.a0(P09D0),
				.a1(P09E0),
				.a2(P09F0),
				.a3(P0AD0),
				.a4(P0AE0),
				.a5(P0AF0),
				.a6(P0BD0),
				.a7(P0BE0),
				.a8(P0BF0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c009D1)
);

ninexnine_unit ninexnine_unit_1006(
				.clk(clk),
				.rstn(rstn),
				.a0(P09D1),
				.a1(P09E1),
				.a2(P09F1),
				.a3(P0AD1),
				.a4(P0AE1),
				.a5(P0AF1),
				.a6(P0BD1),
				.a7(P0BE1),
				.a8(P0BF1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c019D1)
);

ninexnine_unit ninexnine_unit_1007(
				.clk(clk),
				.rstn(rstn),
				.a0(P09D2),
				.a1(P09E2),
				.a2(P09F2),
				.a3(P0AD2),
				.a4(P0AE2),
				.a5(P0AF2),
				.a6(P0BD2),
				.a7(P0BE2),
				.a8(P0BF2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c029D1)
);

assign C09D1=c009D1+c019D1+c029D1;
assign A09D1=(C09D1>=0)?1:0;

ninexnine_unit ninexnine_unit_1008(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A00),
				.a1(P0A10),
				.a2(P0A20),
				.a3(P0B00),
				.a4(P0B10),
				.a5(P0B20),
				.a6(P0C00),
				.a7(P0C10),
				.a8(P0C20),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00A01)
);

ninexnine_unit ninexnine_unit_1009(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A01),
				.a1(P0A11),
				.a2(P0A21),
				.a3(P0B01),
				.a4(P0B11),
				.a5(P0B21),
				.a6(P0C01),
				.a7(P0C11),
				.a8(P0C21),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01A01)
);

ninexnine_unit ninexnine_unit_1010(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A02),
				.a1(P0A12),
				.a2(P0A22),
				.a3(P0B02),
				.a4(P0B12),
				.a5(P0B22),
				.a6(P0C02),
				.a7(P0C12),
				.a8(P0C22),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02A01)
);

assign C0A01=c00A01+c01A01+c02A01;
assign A0A01=(C0A01>=0)?1:0;

ninexnine_unit ninexnine_unit_1011(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A10),
				.a1(P0A20),
				.a2(P0A30),
				.a3(P0B10),
				.a4(P0B20),
				.a5(P0B30),
				.a6(P0C10),
				.a7(P0C20),
				.a8(P0C30),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00A11)
);

ninexnine_unit ninexnine_unit_1012(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A11),
				.a1(P0A21),
				.a2(P0A31),
				.a3(P0B11),
				.a4(P0B21),
				.a5(P0B31),
				.a6(P0C11),
				.a7(P0C21),
				.a8(P0C31),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01A11)
);

ninexnine_unit ninexnine_unit_1013(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A12),
				.a1(P0A22),
				.a2(P0A32),
				.a3(P0B12),
				.a4(P0B22),
				.a5(P0B32),
				.a6(P0C12),
				.a7(P0C22),
				.a8(P0C32),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02A11)
);

assign C0A11=c00A11+c01A11+c02A11;
assign A0A11=(C0A11>=0)?1:0;

ninexnine_unit ninexnine_unit_1014(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A20),
				.a1(P0A30),
				.a2(P0A40),
				.a3(P0B20),
				.a4(P0B30),
				.a5(P0B40),
				.a6(P0C20),
				.a7(P0C30),
				.a8(P0C40),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00A21)
);

ninexnine_unit ninexnine_unit_1015(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A21),
				.a1(P0A31),
				.a2(P0A41),
				.a3(P0B21),
				.a4(P0B31),
				.a5(P0B41),
				.a6(P0C21),
				.a7(P0C31),
				.a8(P0C41),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01A21)
);

ninexnine_unit ninexnine_unit_1016(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A22),
				.a1(P0A32),
				.a2(P0A42),
				.a3(P0B22),
				.a4(P0B32),
				.a5(P0B42),
				.a6(P0C22),
				.a7(P0C32),
				.a8(P0C42),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02A21)
);

assign C0A21=c00A21+c01A21+c02A21;
assign A0A21=(C0A21>=0)?1:0;

ninexnine_unit ninexnine_unit_1017(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A30),
				.a1(P0A40),
				.a2(P0A50),
				.a3(P0B30),
				.a4(P0B40),
				.a5(P0B50),
				.a6(P0C30),
				.a7(P0C40),
				.a8(P0C50),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00A31)
);

ninexnine_unit ninexnine_unit_1018(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A31),
				.a1(P0A41),
				.a2(P0A51),
				.a3(P0B31),
				.a4(P0B41),
				.a5(P0B51),
				.a6(P0C31),
				.a7(P0C41),
				.a8(P0C51),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01A31)
);

ninexnine_unit ninexnine_unit_1019(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A32),
				.a1(P0A42),
				.a2(P0A52),
				.a3(P0B32),
				.a4(P0B42),
				.a5(P0B52),
				.a6(P0C32),
				.a7(P0C42),
				.a8(P0C52),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02A31)
);

assign C0A31=c00A31+c01A31+c02A31;
assign A0A31=(C0A31>=0)?1:0;

ninexnine_unit ninexnine_unit_1020(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A40),
				.a1(P0A50),
				.a2(P0A60),
				.a3(P0B40),
				.a4(P0B50),
				.a5(P0B60),
				.a6(P0C40),
				.a7(P0C50),
				.a8(P0C60),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00A41)
);

ninexnine_unit ninexnine_unit_1021(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A41),
				.a1(P0A51),
				.a2(P0A61),
				.a3(P0B41),
				.a4(P0B51),
				.a5(P0B61),
				.a6(P0C41),
				.a7(P0C51),
				.a8(P0C61),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01A41)
);

ninexnine_unit ninexnine_unit_1022(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A42),
				.a1(P0A52),
				.a2(P0A62),
				.a3(P0B42),
				.a4(P0B52),
				.a5(P0B62),
				.a6(P0C42),
				.a7(P0C52),
				.a8(P0C62),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02A41)
);

assign C0A41=c00A41+c01A41+c02A41;
assign A0A41=(C0A41>=0)?1:0;

ninexnine_unit ninexnine_unit_1023(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A50),
				.a1(P0A60),
				.a2(P0A70),
				.a3(P0B50),
				.a4(P0B60),
				.a5(P0B70),
				.a6(P0C50),
				.a7(P0C60),
				.a8(P0C70),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00A51)
);

ninexnine_unit ninexnine_unit_1024(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A51),
				.a1(P0A61),
				.a2(P0A71),
				.a3(P0B51),
				.a4(P0B61),
				.a5(P0B71),
				.a6(P0C51),
				.a7(P0C61),
				.a8(P0C71),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01A51)
);

ninexnine_unit ninexnine_unit_1025(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A52),
				.a1(P0A62),
				.a2(P0A72),
				.a3(P0B52),
				.a4(P0B62),
				.a5(P0B72),
				.a6(P0C52),
				.a7(P0C62),
				.a8(P0C72),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02A51)
);

assign C0A51=c00A51+c01A51+c02A51;
assign A0A51=(C0A51>=0)?1:0;

ninexnine_unit ninexnine_unit_1026(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A60),
				.a1(P0A70),
				.a2(P0A80),
				.a3(P0B60),
				.a4(P0B70),
				.a5(P0B80),
				.a6(P0C60),
				.a7(P0C70),
				.a8(P0C80),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00A61)
);

ninexnine_unit ninexnine_unit_1027(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A61),
				.a1(P0A71),
				.a2(P0A81),
				.a3(P0B61),
				.a4(P0B71),
				.a5(P0B81),
				.a6(P0C61),
				.a7(P0C71),
				.a8(P0C81),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01A61)
);

ninexnine_unit ninexnine_unit_1028(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A62),
				.a1(P0A72),
				.a2(P0A82),
				.a3(P0B62),
				.a4(P0B72),
				.a5(P0B82),
				.a6(P0C62),
				.a7(P0C72),
				.a8(P0C82),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02A61)
);

assign C0A61=c00A61+c01A61+c02A61;
assign A0A61=(C0A61>=0)?1:0;

ninexnine_unit ninexnine_unit_1029(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A70),
				.a1(P0A80),
				.a2(P0A90),
				.a3(P0B70),
				.a4(P0B80),
				.a5(P0B90),
				.a6(P0C70),
				.a7(P0C80),
				.a8(P0C90),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00A71)
);

ninexnine_unit ninexnine_unit_1030(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A71),
				.a1(P0A81),
				.a2(P0A91),
				.a3(P0B71),
				.a4(P0B81),
				.a5(P0B91),
				.a6(P0C71),
				.a7(P0C81),
				.a8(P0C91),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01A71)
);

ninexnine_unit ninexnine_unit_1031(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A72),
				.a1(P0A82),
				.a2(P0A92),
				.a3(P0B72),
				.a4(P0B82),
				.a5(P0B92),
				.a6(P0C72),
				.a7(P0C82),
				.a8(P0C92),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02A71)
);

assign C0A71=c00A71+c01A71+c02A71;
assign A0A71=(C0A71>=0)?1:0;

ninexnine_unit ninexnine_unit_1032(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A80),
				.a1(P0A90),
				.a2(P0AA0),
				.a3(P0B80),
				.a4(P0B90),
				.a5(P0BA0),
				.a6(P0C80),
				.a7(P0C90),
				.a8(P0CA0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00A81)
);

ninexnine_unit ninexnine_unit_1033(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A81),
				.a1(P0A91),
				.a2(P0AA1),
				.a3(P0B81),
				.a4(P0B91),
				.a5(P0BA1),
				.a6(P0C81),
				.a7(P0C91),
				.a8(P0CA1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01A81)
);

ninexnine_unit ninexnine_unit_1034(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A82),
				.a1(P0A92),
				.a2(P0AA2),
				.a3(P0B82),
				.a4(P0B92),
				.a5(P0BA2),
				.a6(P0C82),
				.a7(P0C92),
				.a8(P0CA2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02A81)
);

assign C0A81=c00A81+c01A81+c02A81;
assign A0A81=(C0A81>=0)?1:0;

ninexnine_unit ninexnine_unit_1035(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A90),
				.a1(P0AA0),
				.a2(P0AB0),
				.a3(P0B90),
				.a4(P0BA0),
				.a5(P0BB0),
				.a6(P0C90),
				.a7(P0CA0),
				.a8(P0CB0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00A91)
);

ninexnine_unit ninexnine_unit_1036(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A91),
				.a1(P0AA1),
				.a2(P0AB1),
				.a3(P0B91),
				.a4(P0BA1),
				.a5(P0BB1),
				.a6(P0C91),
				.a7(P0CA1),
				.a8(P0CB1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01A91)
);

ninexnine_unit ninexnine_unit_1037(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A92),
				.a1(P0AA2),
				.a2(P0AB2),
				.a3(P0B92),
				.a4(P0BA2),
				.a5(P0BB2),
				.a6(P0C92),
				.a7(P0CA2),
				.a8(P0CB2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02A91)
);

assign C0A91=c00A91+c01A91+c02A91;
assign A0A91=(C0A91>=0)?1:0;

ninexnine_unit ninexnine_unit_1038(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AA0),
				.a1(P0AB0),
				.a2(P0AC0),
				.a3(P0BA0),
				.a4(P0BB0),
				.a5(P0BC0),
				.a6(P0CA0),
				.a7(P0CB0),
				.a8(P0CC0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00AA1)
);

ninexnine_unit ninexnine_unit_1039(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AA1),
				.a1(P0AB1),
				.a2(P0AC1),
				.a3(P0BA1),
				.a4(P0BB1),
				.a5(P0BC1),
				.a6(P0CA1),
				.a7(P0CB1),
				.a8(P0CC1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01AA1)
);

ninexnine_unit ninexnine_unit_1040(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AA2),
				.a1(P0AB2),
				.a2(P0AC2),
				.a3(P0BA2),
				.a4(P0BB2),
				.a5(P0BC2),
				.a6(P0CA2),
				.a7(P0CB2),
				.a8(P0CC2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02AA1)
);

assign C0AA1=c00AA1+c01AA1+c02AA1;
assign A0AA1=(C0AA1>=0)?1:0;

ninexnine_unit ninexnine_unit_1041(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AB0),
				.a1(P0AC0),
				.a2(P0AD0),
				.a3(P0BB0),
				.a4(P0BC0),
				.a5(P0BD0),
				.a6(P0CB0),
				.a7(P0CC0),
				.a8(P0CD0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00AB1)
);

ninexnine_unit ninexnine_unit_1042(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AB1),
				.a1(P0AC1),
				.a2(P0AD1),
				.a3(P0BB1),
				.a4(P0BC1),
				.a5(P0BD1),
				.a6(P0CB1),
				.a7(P0CC1),
				.a8(P0CD1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01AB1)
);

ninexnine_unit ninexnine_unit_1043(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AB2),
				.a1(P0AC2),
				.a2(P0AD2),
				.a3(P0BB2),
				.a4(P0BC2),
				.a5(P0BD2),
				.a6(P0CB2),
				.a7(P0CC2),
				.a8(P0CD2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02AB1)
);

assign C0AB1=c00AB1+c01AB1+c02AB1;
assign A0AB1=(C0AB1>=0)?1:0;

ninexnine_unit ninexnine_unit_1044(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AC0),
				.a1(P0AD0),
				.a2(P0AE0),
				.a3(P0BC0),
				.a4(P0BD0),
				.a5(P0BE0),
				.a6(P0CC0),
				.a7(P0CD0),
				.a8(P0CE0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00AC1)
);

ninexnine_unit ninexnine_unit_1045(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AC1),
				.a1(P0AD1),
				.a2(P0AE1),
				.a3(P0BC1),
				.a4(P0BD1),
				.a5(P0BE1),
				.a6(P0CC1),
				.a7(P0CD1),
				.a8(P0CE1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01AC1)
);

ninexnine_unit ninexnine_unit_1046(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AC2),
				.a1(P0AD2),
				.a2(P0AE2),
				.a3(P0BC2),
				.a4(P0BD2),
				.a5(P0BE2),
				.a6(P0CC2),
				.a7(P0CD2),
				.a8(P0CE2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02AC1)
);

assign C0AC1=c00AC1+c01AC1+c02AC1;
assign A0AC1=(C0AC1>=0)?1:0;

ninexnine_unit ninexnine_unit_1047(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AD0),
				.a1(P0AE0),
				.a2(P0AF0),
				.a3(P0BD0),
				.a4(P0BE0),
				.a5(P0BF0),
				.a6(P0CD0),
				.a7(P0CE0),
				.a8(P0CF0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00AD1)
);

ninexnine_unit ninexnine_unit_1048(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AD1),
				.a1(P0AE1),
				.a2(P0AF1),
				.a3(P0BD1),
				.a4(P0BE1),
				.a5(P0BF1),
				.a6(P0CD1),
				.a7(P0CE1),
				.a8(P0CF1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01AD1)
);

ninexnine_unit ninexnine_unit_1049(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AD2),
				.a1(P0AE2),
				.a2(P0AF2),
				.a3(P0BD2),
				.a4(P0BE2),
				.a5(P0BF2),
				.a6(P0CD2),
				.a7(P0CE2),
				.a8(P0CF2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02AD1)
);

assign C0AD1=c00AD1+c01AD1+c02AD1;
assign A0AD1=(C0AD1>=0)?1:0;

ninexnine_unit ninexnine_unit_1050(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B00),
				.a1(P0B10),
				.a2(P0B20),
				.a3(P0C00),
				.a4(P0C10),
				.a5(P0C20),
				.a6(P0D00),
				.a7(P0D10),
				.a8(P0D20),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00B01)
);

ninexnine_unit ninexnine_unit_1051(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B01),
				.a1(P0B11),
				.a2(P0B21),
				.a3(P0C01),
				.a4(P0C11),
				.a5(P0C21),
				.a6(P0D01),
				.a7(P0D11),
				.a8(P0D21),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01B01)
);

ninexnine_unit ninexnine_unit_1052(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B02),
				.a1(P0B12),
				.a2(P0B22),
				.a3(P0C02),
				.a4(P0C12),
				.a5(P0C22),
				.a6(P0D02),
				.a7(P0D12),
				.a8(P0D22),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02B01)
);

assign C0B01=c00B01+c01B01+c02B01;
assign A0B01=(C0B01>=0)?1:0;

ninexnine_unit ninexnine_unit_1053(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B10),
				.a1(P0B20),
				.a2(P0B30),
				.a3(P0C10),
				.a4(P0C20),
				.a5(P0C30),
				.a6(P0D10),
				.a7(P0D20),
				.a8(P0D30),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00B11)
);

ninexnine_unit ninexnine_unit_1054(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B11),
				.a1(P0B21),
				.a2(P0B31),
				.a3(P0C11),
				.a4(P0C21),
				.a5(P0C31),
				.a6(P0D11),
				.a7(P0D21),
				.a8(P0D31),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01B11)
);

ninexnine_unit ninexnine_unit_1055(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B12),
				.a1(P0B22),
				.a2(P0B32),
				.a3(P0C12),
				.a4(P0C22),
				.a5(P0C32),
				.a6(P0D12),
				.a7(P0D22),
				.a8(P0D32),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02B11)
);

assign C0B11=c00B11+c01B11+c02B11;
assign A0B11=(C0B11>=0)?1:0;

ninexnine_unit ninexnine_unit_1056(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B20),
				.a1(P0B30),
				.a2(P0B40),
				.a3(P0C20),
				.a4(P0C30),
				.a5(P0C40),
				.a6(P0D20),
				.a7(P0D30),
				.a8(P0D40),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00B21)
);

ninexnine_unit ninexnine_unit_1057(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B21),
				.a1(P0B31),
				.a2(P0B41),
				.a3(P0C21),
				.a4(P0C31),
				.a5(P0C41),
				.a6(P0D21),
				.a7(P0D31),
				.a8(P0D41),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01B21)
);

ninexnine_unit ninexnine_unit_1058(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B22),
				.a1(P0B32),
				.a2(P0B42),
				.a3(P0C22),
				.a4(P0C32),
				.a5(P0C42),
				.a6(P0D22),
				.a7(P0D32),
				.a8(P0D42),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02B21)
);

assign C0B21=c00B21+c01B21+c02B21;
assign A0B21=(C0B21>=0)?1:0;

ninexnine_unit ninexnine_unit_1059(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B30),
				.a1(P0B40),
				.a2(P0B50),
				.a3(P0C30),
				.a4(P0C40),
				.a5(P0C50),
				.a6(P0D30),
				.a7(P0D40),
				.a8(P0D50),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00B31)
);

ninexnine_unit ninexnine_unit_1060(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B31),
				.a1(P0B41),
				.a2(P0B51),
				.a3(P0C31),
				.a4(P0C41),
				.a5(P0C51),
				.a6(P0D31),
				.a7(P0D41),
				.a8(P0D51),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01B31)
);

ninexnine_unit ninexnine_unit_1061(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B32),
				.a1(P0B42),
				.a2(P0B52),
				.a3(P0C32),
				.a4(P0C42),
				.a5(P0C52),
				.a6(P0D32),
				.a7(P0D42),
				.a8(P0D52),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02B31)
);

assign C0B31=c00B31+c01B31+c02B31;
assign A0B31=(C0B31>=0)?1:0;

ninexnine_unit ninexnine_unit_1062(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B40),
				.a1(P0B50),
				.a2(P0B60),
				.a3(P0C40),
				.a4(P0C50),
				.a5(P0C60),
				.a6(P0D40),
				.a7(P0D50),
				.a8(P0D60),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00B41)
);

ninexnine_unit ninexnine_unit_1063(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B41),
				.a1(P0B51),
				.a2(P0B61),
				.a3(P0C41),
				.a4(P0C51),
				.a5(P0C61),
				.a6(P0D41),
				.a7(P0D51),
				.a8(P0D61),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01B41)
);

ninexnine_unit ninexnine_unit_1064(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B42),
				.a1(P0B52),
				.a2(P0B62),
				.a3(P0C42),
				.a4(P0C52),
				.a5(P0C62),
				.a6(P0D42),
				.a7(P0D52),
				.a8(P0D62),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02B41)
);

assign C0B41=c00B41+c01B41+c02B41;
assign A0B41=(C0B41>=0)?1:0;

ninexnine_unit ninexnine_unit_1065(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B50),
				.a1(P0B60),
				.a2(P0B70),
				.a3(P0C50),
				.a4(P0C60),
				.a5(P0C70),
				.a6(P0D50),
				.a7(P0D60),
				.a8(P0D70),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00B51)
);

ninexnine_unit ninexnine_unit_1066(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B51),
				.a1(P0B61),
				.a2(P0B71),
				.a3(P0C51),
				.a4(P0C61),
				.a5(P0C71),
				.a6(P0D51),
				.a7(P0D61),
				.a8(P0D71),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01B51)
);

ninexnine_unit ninexnine_unit_1067(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B52),
				.a1(P0B62),
				.a2(P0B72),
				.a3(P0C52),
				.a4(P0C62),
				.a5(P0C72),
				.a6(P0D52),
				.a7(P0D62),
				.a8(P0D72),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02B51)
);

assign C0B51=c00B51+c01B51+c02B51;
assign A0B51=(C0B51>=0)?1:0;

ninexnine_unit ninexnine_unit_1068(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B60),
				.a1(P0B70),
				.a2(P0B80),
				.a3(P0C60),
				.a4(P0C70),
				.a5(P0C80),
				.a6(P0D60),
				.a7(P0D70),
				.a8(P0D80),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00B61)
);

ninexnine_unit ninexnine_unit_1069(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B61),
				.a1(P0B71),
				.a2(P0B81),
				.a3(P0C61),
				.a4(P0C71),
				.a5(P0C81),
				.a6(P0D61),
				.a7(P0D71),
				.a8(P0D81),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01B61)
);

ninexnine_unit ninexnine_unit_1070(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B62),
				.a1(P0B72),
				.a2(P0B82),
				.a3(P0C62),
				.a4(P0C72),
				.a5(P0C82),
				.a6(P0D62),
				.a7(P0D72),
				.a8(P0D82),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02B61)
);

assign C0B61=c00B61+c01B61+c02B61;
assign A0B61=(C0B61>=0)?1:0;

ninexnine_unit ninexnine_unit_1071(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B70),
				.a1(P0B80),
				.a2(P0B90),
				.a3(P0C70),
				.a4(P0C80),
				.a5(P0C90),
				.a6(P0D70),
				.a7(P0D80),
				.a8(P0D90),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00B71)
);

ninexnine_unit ninexnine_unit_1072(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B71),
				.a1(P0B81),
				.a2(P0B91),
				.a3(P0C71),
				.a4(P0C81),
				.a5(P0C91),
				.a6(P0D71),
				.a7(P0D81),
				.a8(P0D91),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01B71)
);

ninexnine_unit ninexnine_unit_1073(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B72),
				.a1(P0B82),
				.a2(P0B92),
				.a3(P0C72),
				.a4(P0C82),
				.a5(P0C92),
				.a6(P0D72),
				.a7(P0D82),
				.a8(P0D92),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02B71)
);

assign C0B71=c00B71+c01B71+c02B71;
assign A0B71=(C0B71>=0)?1:0;

ninexnine_unit ninexnine_unit_1074(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B80),
				.a1(P0B90),
				.a2(P0BA0),
				.a3(P0C80),
				.a4(P0C90),
				.a5(P0CA0),
				.a6(P0D80),
				.a7(P0D90),
				.a8(P0DA0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00B81)
);

ninexnine_unit ninexnine_unit_1075(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B81),
				.a1(P0B91),
				.a2(P0BA1),
				.a3(P0C81),
				.a4(P0C91),
				.a5(P0CA1),
				.a6(P0D81),
				.a7(P0D91),
				.a8(P0DA1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01B81)
);

ninexnine_unit ninexnine_unit_1076(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B82),
				.a1(P0B92),
				.a2(P0BA2),
				.a3(P0C82),
				.a4(P0C92),
				.a5(P0CA2),
				.a6(P0D82),
				.a7(P0D92),
				.a8(P0DA2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02B81)
);

assign C0B81=c00B81+c01B81+c02B81;
assign A0B81=(C0B81>=0)?1:0;

ninexnine_unit ninexnine_unit_1077(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B90),
				.a1(P0BA0),
				.a2(P0BB0),
				.a3(P0C90),
				.a4(P0CA0),
				.a5(P0CB0),
				.a6(P0D90),
				.a7(P0DA0),
				.a8(P0DB0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00B91)
);

ninexnine_unit ninexnine_unit_1078(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B91),
				.a1(P0BA1),
				.a2(P0BB1),
				.a3(P0C91),
				.a4(P0CA1),
				.a5(P0CB1),
				.a6(P0D91),
				.a7(P0DA1),
				.a8(P0DB1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01B91)
);

ninexnine_unit ninexnine_unit_1079(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B92),
				.a1(P0BA2),
				.a2(P0BB2),
				.a3(P0C92),
				.a4(P0CA2),
				.a5(P0CB2),
				.a6(P0D92),
				.a7(P0DA2),
				.a8(P0DB2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02B91)
);

assign C0B91=c00B91+c01B91+c02B91;
assign A0B91=(C0B91>=0)?1:0;

ninexnine_unit ninexnine_unit_1080(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BA0),
				.a1(P0BB0),
				.a2(P0BC0),
				.a3(P0CA0),
				.a4(P0CB0),
				.a5(P0CC0),
				.a6(P0DA0),
				.a7(P0DB0),
				.a8(P0DC0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00BA1)
);

ninexnine_unit ninexnine_unit_1081(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BA1),
				.a1(P0BB1),
				.a2(P0BC1),
				.a3(P0CA1),
				.a4(P0CB1),
				.a5(P0CC1),
				.a6(P0DA1),
				.a7(P0DB1),
				.a8(P0DC1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01BA1)
);

ninexnine_unit ninexnine_unit_1082(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BA2),
				.a1(P0BB2),
				.a2(P0BC2),
				.a3(P0CA2),
				.a4(P0CB2),
				.a5(P0CC2),
				.a6(P0DA2),
				.a7(P0DB2),
				.a8(P0DC2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02BA1)
);

assign C0BA1=c00BA1+c01BA1+c02BA1;
assign A0BA1=(C0BA1>=0)?1:0;

ninexnine_unit ninexnine_unit_1083(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BB0),
				.a1(P0BC0),
				.a2(P0BD0),
				.a3(P0CB0),
				.a4(P0CC0),
				.a5(P0CD0),
				.a6(P0DB0),
				.a7(P0DC0),
				.a8(P0DD0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00BB1)
);

ninexnine_unit ninexnine_unit_1084(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BB1),
				.a1(P0BC1),
				.a2(P0BD1),
				.a3(P0CB1),
				.a4(P0CC1),
				.a5(P0CD1),
				.a6(P0DB1),
				.a7(P0DC1),
				.a8(P0DD1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01BB1)
);

ninexnine_unit ninexnine_unit_1085(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BB2),
				.a1(P0BC2),
				.a2(P0BD2),
				.a3(P0CB2),
				.a4(P0CC2),
				.a5(P0CD2),
				.a6(P0DB2),
				.a7(P0DC2),
				.a8(P0DD2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02BB1)
);

assign C0BB1=c00BB1+c01BB1+c02BB1;
assign A0BB1=(C0BB1>=0)?1:0;

ninexnine_unit ninexnine_unit_1086(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BC0),
				.a1(P0BD0),
				.a2(P0BE0),
				.a3(P0CC0),
				.a4(P0CD0),
				.a5(P0CE0),
				.a6(P0DC0),
				.a7(P0DD0),
				.a8(P0DE0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00BC1)
);

ninexnine_unit ninexnine_unit_1087(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BC1),
				.a1(P0BD1),
				.a2(P0BE1),
				.a3(P0CC1),
				.a4(P0CD1),
				.a5(P0CE1),
				.a6(P0DC1),
				.a7(P0DD1),
				.a8(P0DE1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01BC1)
);

ninexnine_unit ninexnine_unit_1088(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BC2),
				.a1(P0BD2),
				.a2(P0BE2),
				.a3(P0CC2),
				.a4(P0CD2),
				.a5(P0CE2),
				.a6(P0DC2),
				.a7(P0DD2),
				.a8(P0DE2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02BC1)
);

assign C0BC1=c00BC1+c01BC1+c02BC1;
assign A0BC1=(C0BC1>=0)?1:0;

ninexnine_unit ninexnine_unit_1089(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BD0),
				.a1(P0BE0),
				.a2(P0BF0),
				.a3(P0CD0),
				.a4(P0CE0),
				.a5(P0CF0),
				.a6(P0DD0),
				.a7(P0DE0),
				.a8(P0DF0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00BD1)
);

ninexnine_unit ninexnine_unit_1090(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BD1),
				.a1(P0BE1),
				.a2(P0BF1),
				.a3(P0CD1),
				.a4(P0CE1),
				.a5(P0CF1),
				.a6(P0DD1),
				.a7(P0DE1),
				.a8(P0DF1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01BD1)
);

ninexnine_unit ninexnine_unit_1091(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BD2),
				.a1(P0BE2),
				.a2(P0BF2),
				.a3(P0CD2),
				.a4(P0CE2),
				.a5(P0CF2),
				.a6(P0DD2),
				.a7(P0DE2),
				.a8(P0DF2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02BD1)
);

assign C0BD1=c00BD1+c01BD1+c02BD1;
assign A0BD1=(C0BD1>=0)?1:0;

ninexnine_unit ninexnine_unit_1092(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C00),
				.a1(P0C10),
				.a2(P0C20),
				.a3(P0D00),
				.a4(P0D10),
				.a5(P0D20),
				.a6(P0E00),
				.a7(P0E10),
				.a8(P0E20),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00C01)
);

ninexnine_unit ninexnine_unit_1093(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C01),
				.a1(P0C11),
				.a2(P0C21),
				.a3(P0D01),
				.a4(P0D11),
				.a5(P0D21),
				.a6(P0E01),
				.a7(P0E11),
				.a8(P0E21),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01C01)
);

ninexnine_unit ninexnine_unit_1094(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C02),
				.a1(P0C12),
				.a2(P0C22),
				.a3(P0D02),
				.a4(P0D12),
				.a5(P0D22),
				.a6(P0E02),
				.a7(P0E12),
				.a8(P0E22),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02C01)
);

assign C0C01=c00C01+c01C01+c02C01;
assign A0C01=(C0C01>=0)?1:0;

ninexnine_unit ninexnine_unit_1095(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C10),
				.a1(P0C20),
				.a2(P0C30),
				.a3(P0D10),
				.a4(P0D20),
				.a5(P0D30),
				.a6(P0E10),
				.a7(P0E20),
				.a8(P0E30),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00C11)
);

ninexnine_unit ninexnine_unit_1096(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C11),
				.a1(P0C21),
				.a2(P0C31),
				.a3(P0D11),
				.a4(P0D21),
				.a5(P0D31),
				.a6(P0E11),
				.a7(P0E21),
				.a8(P0E31),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01C11)
);

ninexnine_unit ninexnine_unit_1097(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C12),
				.a1(P0C22),
				.a2(P0C32),
				.a3(P0D12),
				.a4(P0D22),
				.a5(P0D32),
				.a6(P0E12),
				.a7(P0E22),
				.a8(P0E32),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02C11)
);

assign C0C11=c00C11+c01C11+c02C11;
assign A0C11=(C0C11>=0)?1:0;

ninexnine_unit ninexnine_unit_1098(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C20),
				.a1(P0C30),
				.a2(P0C40),
				.a3(P0D20),
				.a4(P0D30),
				.a5(P0D40),
				.a6(P0E20),
				.a7(P0E30),
				.a8(P0E40),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00C21)
);

ninexnine_unit ninexnine_unit_1099(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C21),
				.a1(P0C31),
				.a2(P0C41),
				.a3(P0D21),
				.a4(P0D31),
				.a5(P0D41),
				.a6(P0E21),
				.a7(P0E31),
				.a8(P0E41),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01C21)
);

ninexnine_unit ninexnine_unit_1100(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C22),
				.a1(P0C32),
				.a2(P0C42),
				.a3(P0D22),
				.a4(P0D32),
				.a5(P0D42),
				.a6(P0E22),
				.a7(P0E32),
				.a8(P0E42),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02C21)
);

assign C0C21=c00C21+c01C21+c02C21;
assign A0C21=(C0C21>=0)?1:0;

ninexnine_unit ninexnine_unit_1101(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C30),
				.a1(P0C40),
				.a2(P0C50),
				.a3(P0D30),
				.a4(P0D40),
				.a5(P0D50),
				.a6(P0E30),
				.a7(P0E40),
				.a8(P0E50),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00C31)
);

ninexnine_unit ninexnine_unit_1102(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C31),
				.a1(P0C41),
				.a2(P0C51),
				.a3(P0D31),
				.a4(P0D41),
				.a5(P0D51),
				.a6(P0E31),
				.a7(P0E41),
				.a8(P0E51),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01C31)
);

ninexnine_unit ninexnine_unit_1103(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C32),
				.a1(P0C42),
				.a2(P0C52),
				.a3(P0D32),
				.a4(P0D42),
				.a5(P0D52),
				.a6(P0E32),
				.a7(P0E42),
				.a8(P0E52),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02C31)
);

assign C0C31=c00C31+c01C31+c02C31;
assign A0C31=(C0C31>=0)?1:0;

ninexnine_unit ninexnine_unit_1104(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C40),
				.a1(P0C50),
				.a2(P0C60),
				.a3(P0D40),
				.a4(P0D50),
				.a5(P0D60),
				.a6(P0E40),
				.a7(P0E50),
				.a8(P0E60),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00C41)
);

ninexnine_unit ninexnine_unit_1105(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C41),
				.a1(P0C51),
				.a2(P0C61),
				.a3(P0D41),
				.a4(P0D51),
				.a5(P0D61),
				.a6(P0E41),
				.a7(P0E51),
				.a8(P0E61),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01C41)
);

ninexnine_unit ninexnine_unit_1106(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C42),
				.a1(P0C52),
				.a2(P0C62),
				.a3(P0D42),
				.a4(P0D52),
				.a5(P0D62),
				.a6(P0E42),
				.a7(P0E52),
				.a8(P0E62),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02C41)
);

assign C0C41=c00C41+c01C41+c02C41;
assign A0C41=(C0C41>=0)?1:0;

ninexnine_unit ninexnine_unit_1107(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C50),
				.a1(P0C60),
				.a2(P0C70),
				.a3(P0D50),
				.a4(P0D60),
				.a5(P0D70),
				.a6(P0E50),
				.a7(P0E60),
				.a8(P0E70),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00C51)
);

ninexnine_unit ninexnine_unit_1108(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C51),
				.a1(P0C61),
				.a2(P0C71),
				.a3(P0D51),
				.a4(P0D61),
				.a5(P0D71),
				.a6(P0E51),
				.a7(P0E61),
				.a8(P0E71),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01C51)
);

ninexnine_unit ninexnine_unit_1109(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C52),
				.a1(P0C62),
				.a2(P0C72),
				.a3(P0D52),
				.a4(P0D62),
				.a5(P0D72),
				.a6(P0E52),
				.a7(P0E62),
				.a8(P0E72),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02C51)
);

assign C0C51=c00C51+c01C51+c02C51;
assign A0C51=(C0C51>=0)?1:0;

ninexnine_unit ninexnine_unit_1110(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C60),
				.a1(P0C70),
				.a2(P0C80),
				.a3(P0D60),
				.a4(P0D70),
				.a5(P0D80),
				.a6(P0E60),
				.a7(P0E70),
				.a8(P0E80),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00C61)
);

ninexnine_unit ninexnine_unit_1111(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C61),
				.a1(P0C71),
				.a2(P0C81),
				.a3(P0D61),
				.a4(P0D71),
				.a5(P0D81),
				.a6(P0E61),
				.a7(P0E71),
				.a8(P0E81),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01C61)
);

ninexnine_unit ninexnine_unit_1112(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C62),
				.a1(P0C72),
				.a2(P0C82),
				.a3(P0D62),
				.a4(P0D72),
				.a5(P0D82),
				.a6(P0E62),
				.a7(P0E72),
				.a8(P0E82),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02C61)
);

assign C0C61=c00C61+c01C61+c02C61;
assign A0C61=(C0C61>=0)?1:0;

ninexnine_unit ninexnine_unit_1113(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C70),
				.a1(P0C80),
				.a2(P0C90),
				.a3(P0D70),
				.a4(P0D80),
				.a5(P0D90),
				.a6(P0E70),
				.a7(P0E80),
				.a8(P0E90),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00C71)
);

ninexnine_unit ninexnine_unit_1114(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C71),
				.a1(P0C81),
				.a2(P0C91),
				.a3(P0D71),
				.a4(P0D81),
				.a5(P0D91),
				.a6(P0E71),
				.a7(P0E81),
				.a8(P0E91),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01C71)
);

ninexnine_unit ninexnine_unit_1115(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C72),
				.a1(P0C82),
				.a2(P0C92),
				.a3(P0D72),
				.a4(P0D82),
				.a5(P0D92),
				.a6(P0E72),
				.a7(P0E82),
				.a8(P0E92),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02C71)
);

assign C0C71=c00C71+c01C71+c02C71;
assign A0C71=(C0C71>=0)?1:0;

ninexnine_unit ninexnine_unit_1116(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C80),
				.a1(P0C90),
				.a2(P0CA0),
				.a3(P0D80),
				.a4(P0D90),
				.a5(P0DA0),
				.a6(P0E80),
				.a7(P0E90),
				.a8(P0EA0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00C81)
);

ninexnine_unit ninexnine_unit_1117(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C81),
				.a1(P0C91),
				.a2(P0CA1),
				.a3(P0D81),
				.a4(P0D91),
				.a5(P0DA1),
				.a6(P0E81),
				.a7(P0E91),
				.a8(P0EA1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01C81)
);

ninexnine_unit ninexnine_unit_1118(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C82),
				.a1(P0C92),
				.a2(P0CA2),
				.a3(P0D82),
				.a4(P0D92),
				.a5(P0DA2),
				.a6(P0E82),
				.a7(P0E92),
				.a8(P0EA2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02C81)
);

assign C0C81=c00C81+c01C81+c02C81;
assign A0C81=(C0C81>=0)?1:0;

ninexnine_unit ninexnine_unit_1119(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C90),
				.a1(P0CA0),
				.a2(P0CB0),
				.a3(P0D90),
				.a4(P0DA0),
				.a5(P0DB0),
				.a6(P0E90),
				.a7(P0EA0),
				.a8(P0EB0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00C91)
);

ninexnine_unit ninexnine_unit_1120(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C91),
				.a1(P0CA1),
				.a2(P0CB1),
				.a3(P0D91),
				.a4(P0DA1),
				.a5(P0DB1),
				.a6(P0E91),
				.a7(P0EA1),
				.a8(P0EB1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01C91)
);

ninexnine_unit ninexnine_unit_1121(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C92),
				.a1(P0CA2),
				.a2(P0CB2),
				.a3(P0D92),
				.a4(P0DA2),
				.a5(P0DB2),
				.a6(P0E92),
				.a7(P0EA2),
				.a8(P0EB2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02C91)
);

assign C0C91=c00C91+c01C91+c02C91;
assign A0C91=(C0C91>=0)?1:0;

ninexnine_unit ninexnine_unit_1122(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CA0),
				.a1(P0CB0),
				.a2(P0CC0),
				.a3(P0DA0),
				.a4(P0DB0),
				.a5(P0DC0),
				.a6(P0EA0),
				.a7(P0EB0),
				.a8(P0EC0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00CA1)
);

ninexnine_unit ninexnine_unit_1123(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CA1),
				.a1(P0CB1),
				.a2(P0CC1),
				.a3(P0DA1),
				.a4(P0DB1),
				.a5(P0DC1),
				.a6(P0EA1),
				.a7(P0EB1),
				.a8(P0EC1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01CA1)
);

ninexnine_unit ninexnine_unit_1124(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CA2),
				.a1(P0CB2),
				.a2(P0CC2),
				.a3(P0DA2),
				.a4(P0DB2),
				.a5(P0DC2),
				.a6(P0EA2),
				.a7(P0EB2),
				.a8(P0EC2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02CA1)
);

assign C0CA1=c00CA1+c01CA1+c02CA1;
assign A0CA1=(C0CA1>=0)?1:0;

ninexnine_unit ninexnine_unit_1125(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CB0),
				.a1(P0CC0),
				.a2(P0CD0),
				.a3(P0DB0),
				.a4(P0DC0),
				.a5(P0DD0),
				.a6(P0EB0),
				.a7(P0EC0),
				.a8(P0ED0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00CB1)
);

ninexnine_unit ninexnine_unit_1126(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CB1),
				.a1(P0CC1),
				.a2(P0CD1),
				.a3(P0DB1),
				.a4(P0DC1),
				.a5(P0DD1),
				.a6(P0EB1),
				.a7(P0EC1),
				.a8(P0ED1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01CB1)
);

ninexnine_unit ninexnine_unit_1127(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CB2),
				.a1(P0CC2),
				.a2(P0CD2),
				.a3(P0DB2),
				.a4(P0DC2),
				.a5(P0DD2),
				.a6(P0EB2),
				.a7(P0EC2),
				.a8(P0ED2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02CB1)
);

assign C0CB1=c00CB1+c01CB1+c02CB1;
assign A0CB1=(C0CB1>=0)?1:0;

ninexnine_unit ninexnine_unit_1128(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CC0),
				.a1(P0CD0),
				.a2(P0CE0),
				.a3(P0DC0),
				.a4(P0DD0),
				.a5(P0DE0),
				.a6(P0EC0),
				.a7(P0ED0),
				.a8(P0EE0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00CC1)
);

ninexnine_unit ninexnine_unit_1129(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CC1),
				.a1(P0CD1),
				.a2(P0CE1),
				.a3(P0DC1),
				.a4(P0DD1),
				.a5(P0DE1),
				.a6(P0EC1),
				.a7(P0ED1),
				.a8(P0EE1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01CC1)
);

ninexnine_unit ninexnine_unit_1130(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CC2),
				.a1(P0CD2),
				.a2(P0CE2),
				.a3(P0DC2),
				.a4(P0DD2),
				.a5(P0DE2),
				.a6(P0EC2),
				.a7(P0ED2),
				.a8(P0EE2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02CC1)
);

assign C0CC1=c00CC1+c01CC1+c02CC1;
assign A0CC1=(C0CC1>=0)?1:0;

ninexnine_unit ninexnine_unit_1131(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CD0),
				.a1(P0CE0),
				.a2(P0CF0),
				.a3(P0DD0),
				.a4(P0DE0),
				.a5(P0DF0),
				.a6(P0ED0),
				.a7(P0EE0),
				.a8(P0EF0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00CD1)
);

ninexnine_unit ninexnine_unit_1132(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CD1),
				.a1(P0CE1),
				.a2(P0CF1),
				.a3(P0DD1),
				.a4(P0DE1),
				.a5(P0DF1),
				.a6(P0ED1),
				.a7(P0EE1),
				.a8(P0EF1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01CD1)
);

ninexnine_unit ninexnine_unit_1133(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CD2),
				.a1(P0CE2),
				.a2(P0CF2),
				.a3(P0DD2),
				.a4(P0DE2),
				.a5(P0DF2),
				.a6(P0ED2),
				.a7(P0EE2),
				.a8(P0EF2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02CD1)
);

assign C0CD1=c00CD1+c01CD1+c02CD1;
assign A0CD1=(C0CD1>=0)?1:0;

ninexnine_unit ninexnine_unit_1134(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D00),
				.a1(P0D10),
				.a2(P0D20),
				.a3(P0E00),
				.a4(P0E10),
				.a5(P0E20),
				.a6(P0F00),
				.a7(P0F10),
				.a8(P0F20),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00D01)
);

ninexnine_unit ninexnine_unit_1135(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D01),
				.a1(P0D11),
				.a2(P0D21),
				.a3(P0E01),
				.a4(P0E11),
				.a5(P0E21),
				.a6(P0F01),
				.a7(P0F11),
				.a8(P0F21),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01D01)
);

ninexnine_unit ninexnine_unit_1136(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D02),
				.a1(P0D12),
				.a2(P0D22),
				.a3(P0E02),
				.a4(P0E12),
				.a5(P0E22),
				.a6(P0F02),
				.a7(P0F12),
				.a8(P0F22),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02D01)
);

assign C0D01=c00D01+c01D01+c02D01;
assign A0D01=(C0D01>=0)?1:0;

ninexnine_unit ninexnine_unit_1137(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D10),
				.a1(P0D20),
				.a2(P0D30),
				.a3(P0E10),
				.a4(P0E20),
				.a5(P0E30),
				.a6(P0F10),
				.a7(P0F20),
				.a8(P0F30),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00D11)
);

ninexnine_unit ninexnine_unit_1138(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D11),
				.a1(P0D21),
				.a2(P0D31),
				.a3(P0E11),
				.a4(P0E21),
				.a5(P0E31),
				.a6(P0F11),
				.a7(P0F21),
				.a8(P0F31),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01D11)
);

ninexnine_unit ninexnine_unit_1139(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D12),
				.a1(P0D22),
				.a2(P0D32),
				.a3(P0E12),
				.a4(P0E22),
				.a5(P0E32),
				.a6(P0F12),
				.a7(P0F22),
				.a8(P0F32),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02D11)
);

assign C0D11=c00D11+c01D11+c02D11;
assign A0D11=(C0D11>=0)?1:0;

ninexnine_unit ninexnine_unit_1140(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D20),
				.a1(P0D30),
				.a2(P0D40),
				.a3(P0E20),
				.a4(P0E30),
				.a5(P0E40),
				.a6(P0F20),
				.a7(P0F30),
				.a8(P0F40),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00D21)
);

ninexnine_unit ninexnine_unit_1141(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D21),
				.a1(P0D31),
				.a2(P0D41),
				.a3(P0E21),
				.a4(P0E31),
				.a5(P0E41),
				.a6(P0F21),
				.a7(P0F31),
				.a8(P0F41),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01D21)
);

ninexnine_unit ninexnine_unit_1142(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D22),
				.a1(P0D32),
				.a2(P0D42),
				.a3(P0E22),
				.a4(P0E32),
				.a5(P0E42),
				.a6(P0F22),
				.a7(P0F32),
				.a8(P0F42),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02D21)
);

assign C0D21=c00D21+c01D21+c02D21;
assign A0D21=(C0D21>=0)?1:0;

ninexnine_unit ninexnine_unit_1143(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D30),
				.a1(P0D40),
				.a2(P0D50),
				.a3(P0E30),
				.a4(P0E40),
				.a5(P0E50),
				.a6(P0F30),
				.a7(P0F40),
				.a8(P0F50),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00D31)
);

ninexnine_unit ninexnine_unit_1144(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D31),
				.a1(P0D41),
				.a2(P0D51),
				.a3(P0E31),
				.a4(P0E41),
				.a5(P0E51),
				.a6(P0F31),
				.a7(P0F41),
				.a8(P0F51),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01D31)
);

ninexnine_unit ninexnine_unit_1145(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D32),
				.a1(P0D42),
				.a2(P0D52),
				.a3(P0E32),
				.a4(P0E42),
				.a5(P0E52),
				.a6(P0F32),
				.a7(P0F42),
				.a8(P0F52),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02D31)
);

assign C0D31=c00D31+c01D31+c02D31;
assign A0D31=(C0D31>=0)?1:0;

ninexnine_unit ninexnine_unit_1146(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D40),
				.a1(P0D50),
				.a2(P0D60),
				.a3(P0E40),
				.a4(P0E50),
				.a5(P0E60),
				.a6(P0F40),
				.a7(P0F50),
				.a8(P0F60),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00D41)
);

ninexnine_unit ninexnine_unit_1147(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D41),
				.a1(P0D51),
				.a2(P0D61),
				.a3(P0E41),
				.a4(P0E51),
				.a5(P0E61),
				.a6(P0F41),
				.a7(P0F51),
				.a8(P0F61),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01D41)
);

ninexnine_unit ninexnine_unit_1148(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D42),
				.a1(P0D52),
				.a2(P0D62),
				.a3(P0E42),
				.a4(P0E52),
				.a5(P0E62),
				.a6(P0F42),
				.a7(P0F52),
				.a8(P0F62),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02D41)
);

assign C0D41=c00D41+c01D41+c02D41;
assign A0D41=(C0D41>=0)?1:0;

ninexnine_unit ninexnine_unit_1149(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D50),
				.a1(P0D60),
				.a2(P0D70),
				.a3(P0E50),
				.a4(P0E60),
				.a5(P0E70),
				.a6(P0F50),
				.a7(P0F60),
				.a8(P0F70),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00D51)
);

ninexnine_unit ninexnine_unit_1150(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D51),
				.a1(P0D61),
				.a2(P0D71),
				.a3(P0E51),
				.a4(P0E61),
				.a5(P0E71),
				.a6(P0F51),
				.a7(P0F61),
				.a8(P0F71),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01D51)
);

ninexnine_unit ninexnine_unit_1151(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D52),
				.a1(P0D62),
				.a2(P0D72),
				.a3(P0E52),
				.a4(P0E62),
				.a5(P0E72),
				.a6(P0F52),
				.a7(P0F62),
				.a8(P0F72),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02D51)
);

assign C0D51=c00D51+c01D51+c02D51;
assign A0D51=(C0D51>=0)?1:0;

ninexnine_unit ninexnine_unit_1152(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D60),
				.a1(P0D70),
				.a2(P0D80),
				.a3(P0E60),
				.a4(P0E70),
				.a5(P0E80),
				.a6(P0F60),
				.a7(P0F70),
				.a8(P0F80),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00D61)
);

ninexnine_unit ninexnine_unit_1153(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D61),
				.a1(P0D71),
				.a2(P0D81),
				.a3(P0E61),
				.a4(P0E71),
				.a5(P0E81),
				.a6(P0F61),
				.a7(P0F71),
				.a8(P0F81),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01D61)
);

ninexnine_unit ninexnine_unit_1154(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D62),
				.a1(P0D72),
				.a2(P0D82),
				.a3(P0E62),
				.a4(P0E72),
				.a5(P0E82),
				.a6(P0F62),
				.a7(P0F72),
				.a8(P0F82),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02D61)
);

assign C0D61=c00D61+c01D61+c02D61;
assign A0D61=(C0D61>=0)?1:0;

ninexnine_unit ninexnine_unit_1155(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D70),
				.a1(P0D80),
				.a2(P0D90),
				.a3(P0E70),
				.a4(P0E80),
				.a5(P0E90),
				.a6(P0F70),
				.a7(P0F80),
				.a8(P0F90),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00D71)
);

ninexnine_unit ninexnine_unit_1156(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D71),
				.a1(P0D81),
				.a2(P0D91),
				.a3(P0E71),
				.a4(P0E81),
				.a5(P0E91),
				.a6(P0F71),
				.a7(P0F81),
				.a8(P0F91),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01D71)
);

ninexnine_unit ninexnine_unit_1157(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D72),
				.a1(P0D82),
				.a2(P0D92),
				.a3(P0E72),
				.a4(P0E82),
				.a5(P0E92),
				.a6(P0F72),
				.a7(P0F82),
				.a8(P0F92),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02D71)
);

assign C0D71=c00D71+c01D71+c02D71;
assign A0D71=(C0D71>=0)?1:0;

ninexnine_unit ninexnine_unit_1158(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D80),
				.a1(P0D90),
				.a2(P0DA0),
				.a3(P0E80),
				.a4(P0E90),
				.a5(P0EA0),
				.a6(P0F80),
				.a7(P0F90),
				.a8(P0FA0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00D81)
);

ninexnine_unit ninexnine_unit_1159(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D81),
				.a1(P0D91),
				.a2(P0DA1),
				.a3(P0E81),
				.a4(P0E91),
				.a5(P0EA1),
				.a6(P0F81),
				.a7(P0F91),
				.a8(P0FA1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01D81)
);

ninexnine_unit ninexnine_unit_1160(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D82),
				.a1(P0D92),
				.a2(P0DA2),
				.a3(P0E82),
				.a4(P0E92),
				.a5(P0EA2),
				.a6(P0F82),
				.a7(P0F92),
				.a8(P0FA2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02D81)
);

assign C0D81=c00D81+c01D81+c02D81;
assign A0D81=(C0D81>=0)?1:0;

ninexnine_unit ninexnine_unit_1161(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D90),
				.a1(P0DA0),
				.a2(P0DB0),
				.a3(P0E90),
				.a4(P0EA0),
				.a5(P0EB0),
				.a6(P0F90),
				.a7(P0FA0),
				.a8(P0FB0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00D91)
);

ninexnine_unit ninexnine_unit_1162(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D91),
				.a1(P0DA1),
				.a2(P0DB1),
				.a3(P0E91),
				.a4(P0EA1),
				.a5(P0EB1),
				.a6(P0F91),
				.a7(P0FA1),
				.a8(P0FB1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01D91)
);

ninexnine_unit ninexnine_unit_1163(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D92),
				.a1(P0DA2),
				.a2(P0DB2),
				.a3(P0E92),
				.a4(P0EA2),
				.a5(P0EB2),
				.a6(P0F92),
				.a7(P0FA2),
				.a8(P0FB2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02D91)
);

assign C0D91=c00D91+c01D91+c02D91;
assign A0D91=(C0D91>=0)?1:0;

ninexnine_unit ninexnine_unit_1164(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DA0),
				.a1(P0DB0),
				.a2(P0DC0),
				.a3(P0EA0),
				.a4(P0EB0),
				.a5(P0EC0),
				.a6(P0FA0),
				.a7(P0FB0),
				.a8(P0FC0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00DA1)
);

ninexnine_unit ninexnine_unit_1165(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DA1),
				.a1(P0DB1),
				.a2(P0DC1),
				.a3(P0EA1),
				.a4(P0EB1),
				.a5(P0EC1),
				.a6(P0FA1),
				.a7(P0FB1),
				.a8(P0FC1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01DA1)
);

ninexnine_unit ninexnine_unit_1166(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DA2),
				.a1(P0DB2),
				.a2(P0DC2),
				.a3(P0EA2),
				.a4(P0EB2),
				.a5(P0EC2),
				.a6(P0FA2),
				.a7(P0FB2),
				.a8(P0FC2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02DA1)
);

assign C0DA1=c00DA1+c01DA1+c02DA1;
assign A0DA1=(C0DA1>=0)?1:0;

ninexnine_unit ninexnine_unit_1167(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DB0),
				.a1(P0DC0),
				.a2(P0DD0),
				.a3(P0EB0),
				.a4(P0EC0),
				.a5(P0ED0),
				.a6(P0FB0),
				.a7(P0FC0),
				.a8(P0FD0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00DB1)
);

ninexnine_unit ninexnine_unit_1168(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DB1),
				.a1(P0DC1),
				.a2(P0DD1),
				.a3(P0EB1),
				.a4(P0EC1),
				.a5(P0ED1),
				.a6(P0FB1),
				.a7(P0FC1),
				.a8(P0FD1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01DB1)
);

ninexnine_unit ninexnine_unit_1169(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DB2),
				.a1(P0DC2),
				.a2(P0DD2),
				.a3(P0EB2),
				.a4(P0EC2),
				.a5(P0ED2),
				.a6(P0FB2),
				.a7(P0FC2),
				.a8(P0FD2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02DB1)
);

assign C0DB1=c00DB1+c01DB1+c02DB1;
assign A0DB1=(C0DB1>=0)?1:0;

ninexnine_unit ninexnine_unit_1170(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DC0),
				.a1(P0DD0),
				.a2(P0DE0),
				.a3(P0EC0),
				.a4(P0ED0),
				.a5(P0EE0),
				.a6(P0FC0),
				.a7(P0FD0),
				.a8(P0FE0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00DC1)
);

ninexnine_unit ninexnine_unit_1171(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DC1),
				.a1(P0DD1),
				.a2(P0DE1),
				.a3(P0EC1),
				.a4(P0ED1),
				.a5(P0EE1),
				.a6(P0FC1),
				.a7(P0FD1),
				.a8(P0FE1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01DC1)
);

ninexnine_unit ninexnine_unit_1172(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DC2),
				.a1(P0DD2),
				.a2(P0DE2),
				.a3(P0EC2),
				.a4(P0ED2),
				.a5(P0EE2),
				.a6(P0FC2),
				.a7(P0FD2),
				.a8(P0FE2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02DC1)
);

assign C0DC1=c00DC1+c01DC1+c02DC1;
assign A0DC1=(C0DC1>=0)?1:0;

ninexnine_unit ninexnine_unit_1173(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DD0),
				.a1(P0DE0),
				.a2(P0DF0),
				.a3(P0ED0),
				.a4(P0EE0),
				.a5(P0EF0),
				.a6(P0FD0),
				.a7(P0FE0),
				.a8(P0FF0),
				.b0(W01000),
				.b1(W01010),
				.b2(W01020),
				.b3(W01100),
				.b4(W01110),
				.b5(W01120),
				.b6(W01200),
				.b7(W01210),
				.b8(W01220),
				.c(c00DD1)
);

ninexnine_unit ninexnine_unit_1174(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DD1),
				.a1(P0DE1),
				.a2(P0DF1),
				.a3(P0ED1),
				.a4(P0EE1),
				.a5(P0EF1),
				.a6(P0FD1),
				.a7(P0FE1),
				.a8(P0FF1),
				.b0(W01001),
				.b1(W01011),
				.b2(W01021),
				.b3(W01101),
				.b4(W01111),
				.b5(W01121),
				.b6(W01201),
				.b7(W01211),
				.b8(W01221),
				.c(c01DD1)
);

ninexnine_unit ninexnine_unit_1175(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DD2),
				.a1(P0DE2),
				.a2(P0DF2),
				.a3(P0ED2),
				.a4(P0EE2),
				.a5(P0EF2),
				.a6(P0FD2),
				.a7(P0FE2),
				.a8(P0FF2),
				.b0(W01002),
				.b1(W01012),
				.b2(W01022),
				.b3(W01102),
				.b4(W01112),
				.b5(W01122),
				.b6(W01202),
				.b7(W01212),
				.b8(W01222),
				.c(c02DD1)
);

assign C0DD1=c00DD1+c01DD1+c02DD1;
assign A0DD1=(C0DD1>=0)?1:0;

ninexnine_unit ninexnine_unit_1176(
				.clk(clk),
				.rstn(rstn),
				.a0(P0000),
				.a1(P0010),
				.a2(P0020),
				.a3(P0100),
				.a4(P0110),
				.a5(P0120),
				.a6(P0200),
				.a7(P0210),
				.a8(P0220),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00002)
);

ninexnine_unit ninexnine_unit_1177(
				.clk(clk),
				.rstn(rstn),
				.a0(P0001),
				.a1(P0011),
				.a2(P0021),
				.a3(P0101),
				.a4(P0111),
				.a5(P0121),
				.a6(P0201),
				.a7(P0211),
				.a8(P0221),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01002)
);

ninexnine_unit ninexnine_unit_1178(
				.clk(clk),
				.rstn(rstn),
				.a0(P0002),
				.a1(P0012),
				.a2(P0022),
				.a3(P0102),
				.a4(P0112),
				.a5(P0122),
				.a6(P0202),
				.a7(P0212),
				.a8(P0222),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02002)
);

assign C0002=c00002+c01002+c02002;
assign A0002=(C0002>=0)?1:0;

ninexnine_unit ninexnine_unit_1179(
				.clk(clk),
				.rstn(rstn),
				.a0(P0010),
				.a1(P0020),
				.a2(P0030),
				.a3(P0110),
				.a4(P0120),
				.a5(P0130),
				.a6(P0210),
				.a7(P0220),
				.a8(P0230),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00012)
);

ninexnine_unit ninexnine_unit_1180(
				.clk(clk),
				.rstn(rstn),
				.a0(P0011),
				.a1(P0021),
				.a2(P0031),
				.a3(P0111),
				.a4(P0121),
				.a5(P0131),
				.a6(P0211),
				.a7(P0221),
				.a8(P0231),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01012)
);

ninexnine_unit ninexnine_unit_1181(
				.clk(clk),
				.rstn(rstn),
				.a0(P0012),
				.a1(P0022),
				.a2(P0032),
				.a3(P0112),
				.a4(P0122),
				.a5(P0132),
				.a6(P0212),
				.a7(P0222),
				.a8(P0232),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02012)
);

assign C0012=c00012+c01012+c02012;
assign A0012=(C0012>=0)?1:0;

ninexnine_unit ninexnine_unit_1182(
				.clk(clk),
				.rstn(rstn),
				.a0(P0020),
				.a1(P0030),
				.a2(P0040),
				.a3(P0120),
				.a4(P0130),
				.a5(P0140),
				.a6(P0220),
				.a7(P0230),
				.a8(P0240),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00022)
);

ninexnine_unit ninexnine_unit_1183(
				.clk(clk),
				.rstn(rstn),
				.a0(P0021),
				.a1(P0031),
				.a2(P0041),
				.a3(P0121),
				.a4(P0131),
				.a5(P0141),
				.a6(P0221),
				.a7(P0231),
				.a8(P0241),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01022)
);

ninexnine_unit ninexnine_unit_1184(
				.clk(clk),
				.rstn(rstn),
				.a0(P0022),
				.a1(P0032),
				.a2(P0042),
				.a3(P0122),
				.a4(P0132),
				.a5(P0142),
				.a6(P0222),
				.a7(P0232),
				.a8(P0242),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02022)
);

assign C0022=c00022+c01022+c02022;
assign A0022=(C0022>=0)?1:0;

ninexnine_unit ninexnine_unit_1185(
				.clk(clk),
				.rstn(rstn),
				.a0(P0030),
				.a1(P0040),
				.a2(P0050),
				.a3(P0130),
				.a4(P0140),
				.a5(P0150),
				.a6(P0230),
				.a7(P0240),
				.a8(P0250),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00032)
);

ninexnine_unit ninexnine_unit_1186(
				.clk(clk),
				.rstn(rstn),
				.a0(P0031),
				.a1(P0041),
				.a2(P0051),
				.a3(P0131),
				.a4(P0141),
				.a5(P0151),
				.a6(P0231),
				.a7(P0241),
				.a8(P0251),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01032)
);

ninexnine_unit ninexnine_unit_1187(
				.clk(clk),
				.rstn(rstn),
				.a0(P0032),
				.a1(P0042),
				.a2(P0052),
				.a3(P0132),
				.a4(P0142),
				.a5(P0152),
				.a6(P0232),
				.a7(P0242),
				.a8(P0252),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02032)
);

assign C0032=c00032+c01032+c02032;
assign A0032=(C0032>=0)?1:0;

ninexnine_unit ninexnine_unit_1188(
				.clk(clk),
				.rstn(rstn),
				.a0(P0040),
				.a1(P0050),
				.a2(P0060),
				.a3(P0140),
				.a4(P0150),
				.a5(P0160),
				.a6(P0240),
				.a7(P0250),
				.a8(P0260),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00042)
);

ninexnine_unit ninexnine_unit_1189(
				.clk(clk),
				.rstn(rstn),
				.a0(P0041),
				.a1(P0051),
				.a2(P0061),
				.a3(P0141),
				.a4(P0151),
				.a5(P0161),
				.a6(P0241),
				.a7(P0251),
				.a8(P0261),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01042)
);

ninexnine_unit ninexnine_unit_1190(
				.clk(clk),
				.rstn(rstn),
				.a0(P0042),
				.a1(P0052),
				.a2(P0062),
				.a3(P0142),
				.a4(P0152),
				.a5(P0162),
				.a6(P0242),
				.a7(P0252),
				.a8(P0262),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02042)
);

assign C0042=c00042+c01042+c02042;
assign A0042=(C0042>=0)?1:0;

ninexnine_unit ninexnine_unit_1191(
				.clk(clk),
				.rstn(rstn),
				.a0(P0050),
				.a1(P0060),
				.a2(P0070),
				.a3(P0150),
				.a4(P0160),
				.a5(P0170),
				.a6(P0250),
				.a7(P0260),
				.a8(P0270),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00052)
);

ninexnine_unit ninexnine_unit_1192(
				.clk(clk),
				.rstn(rstn),
				.a0(P0051),
				.a1(P0061),
				.a2(P0071),
				.a3(P0151),
				.a4(P0161),
				.a5(P0171),
				.a6(P0251),
				.a7(P0261),
				.a8(P0271),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01052)
);

ninexnine_unit ninexnine_unit_1193(
				.clk(clk),
				.rstn(rstn),
				.a0(P0052),
				.a1(P0062),
				.a2(P0072),
				.a3(P0152),
				.a4(P0162),
				.a5(P0172),
				.a6(P0252),
				.a7(P0262),
				.a8(P0272),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02052)
);

assign C0052=c00052+c01052+c02052;
assign A0052=(C0052>=0)?1:0;

ninexnine_unit ninexnine_unit_1194(
				.clk(clk),
				.rstn(rstn),
				.a0(P0060),
				.a1(P0070),
				.a2(P0080),
				.a3(P0160),
				.a4(P0170),
				.a5(P0180),
				.a6(P0260),
				.a7(P0270),
				.a8(P0280),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00062)
);

ninexnine_unit ninexnine_unit_1195(
				.clk(clk),
				.rstn(rstn),
				.a0(P0061),
				.a1(P0071),
				.a2(P0081),
				.a3(P0161),
				.a4(P0171),
				.a5(P0181),
				.a6(P0261),
				.a7(P0271),
				.a8(P0281),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01062)
);

ninexnine_unit ninexnine_unit_1196(
				.clk(clk),
				.rstn(rstn),
				.a0(P0062),
				.a1(P0072),
				.a2(P0082),
				.a3(P0162),
				.a4(P0172),
				.a5(P0182),
				.a6(P0262),
				.a7(P0272),
				.a8(P0282),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02062)
);

assign C0062=c00062+c01062+c02062;
assign A0062=(C0062>=0)?1:0;

ninexnine_unit ninexnine_unit_1197(
				.clk(clk),
				.rstn(rstn),
				.a0(P0070),
				.a1(P0080),
				.a2(P0090),
				.a3(P0170),
				.a4(P0180),
				.a5(P0190),
				.a6(P0270),
				.a7(P0280),
				.a8(P0290),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00072)
);

ninexnine_unit ninexnine_unit_1198(
				.clk(clk),
				.rstn(rstn),
				.a0(P0071),
				.a1(P0081),
				.a2(P0091),
				.a3(P0171),
				.a4(P0181),
				.a5(P0191),
				.a6(P0271),
				.a7(P0281),
				.a8(P0291),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01072)
);

ninexnine_unit ninexnine_unit_1199(
				.clk(clk),
				.rstn(rstn),
				.a0(P0072),
				.a1(P0082),
				.a2(P0092),
				.a3(P0172),
				.a4(P0182),
				.a5(P0192),
				.a6(P0272),
				.a7(P0282),
				.a8(P0292),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02072)
);

assign C0072=c00072+c01072+c02072;
assign A0072=(C0072>=0)?1:0;

ninexnine_unit ninexnine_unit_1200(
				.clk(clk),
				.rstn(rstn),
				.a0(P0080),
				.a1(P0090),
				.a2(P00A0),
				.a3(P0180),
				.a4(P0190),
				.a5(P01A0),
				.a6(P0280),
				.a7(P0290),
				.a8(P02A0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00082)
);

ninexnine_unit ninexnine_unit_1201(
				.clk(clk),
				.rstn(rstn),
				.a0(P0081),
				.a1(P0091),
				.a2(P00A1),
				.a3(P0181),
				.a4(P0191),
				.a5(P01A1),
				.a6(P0281),
				.a7(P0291),
				.a8(P02A1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01082)
);

ninexnine_unit ninexnine_unit_1202(
				.clk(clk),
				.rstn(rstn),
				.a0(P0082),
				.a1(P0092),
				.a2(P00A2),
				.a3(P0182),
				.a4(P0192),
				.a5(P01A2),
				.a6(P0282),
				.a7(P0292),
				.a8(P02A2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02082)
);

assign C0082=c00082+c01082+c02082;
assign A0082=(C0082>=0)?1:0;

ninexnine_unit ninexnine_unit_1203(
				.clk(clk),
				.rstn(rstn),
				.a0(P0090),
				.a1(P00A0),
				.a2(P00B0),
				.a3(P0190),
				.a4(P01A0),
				.a5(P01B0),
				.a6(P0290),
				.a7(P02A0),
				.a8(P02B0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00092)
);

ninexnine_unit ninexnine_unit_1204(
				.clk(clk),
				.rstn(rstn),
				.a0(P0091),
				.a1(P00A1),
				.a2(P00B1),
				.a3(P0191),
				.a4(P01A1),
				.a5(P01B1),
				.a6(P0291),
				.a7(P02A1),
				.a8(P02B1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01092)
);

ninexnine_unit ninexnine_unit_1205(
				.clk(clk),
				.rstn(rstn),
				.a0(P0092),
				.a1(P00A2),
				.a2(P00B2),
				.a3(P0192),
				.a4(P01A2),
				.a5(P01B2),
				.a6(P0292),
				.a7(P02A2),
				.a8(P02B2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02092)
);

assign C0092=c00092+c01092+c02092;
assign A0092=(C0092>=0)?1:0;

ninexnine_unit ninexnine_unit_1206(
				.clk(clk),
				.rstn(rstn),
				.a0(P00A0),
				.a1(P00B0),
				.a2(P00C0),
				.a3(P01A0),
				.a4(P01B0),
				.a5(P01C0),
				.a6(P02A0),
				.a7(P02B0),
				.a8(P02C0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c000A2)
);

ninexnine_unit ninexnine_unit_1207(
				.clk(clk),
				.rstn(rstn),
				.a0(P00A1),
				.a1(P00B1),
				.a2(P00C1),
				.a3(P01A1),
				.a4(P01B1),
				.a5(P01C1),
				.a6(P02A1),
				.a7(P02B1),
				.a8(P02C1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c010A2)
);

ninexnine_unit ninexnine_unit_1208(
				.clk(clk),
				.rstn(rstn),
				.a0(P00A2),
				.a1(P00B2),
				.a2(P00C2),
				.a3(P01A2),
				.a4(P01B2),
				.a5(P01C2),
				.a6(P02A2),
				.a7(P02B2),
				.a8(P02C2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c020A2)
);

assign C00A2=c000A2+c010A2+c020A2;
assign A00A2=(C00A2>=0)?1:0;

ninexnine_unit ninexnine_unit_1209(
				.clk(clk),
				.rstn(rstn),
				.a0(P00B0),
				.a1(P00C0),
				.a2(P00D0),
				.a3(P01B0),
				.a4(P01C0),
				.a5(P01D0),
				.a6(P02B0),
				.a7(P02C0),
				.a8(P02D0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c000B2)
);

ninexnine_unit ninexnine_unit_1210(
				.clk(clk),
				.rstn(rstn),
				.a0(P00B1),
				.a1(P00C1),
				.a2(P00D1),
				.a3(P01B1),
				.a4(P01C1),
				.a5(P01D1),
				.a6(P02B1),
				.a7(P02C1),
				.a8(P02D1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c010B2)
);

ninexnine_unit ninexnine_unit_1211(
				.clk(clk),
				.rstn(rstn),
				.a0(P00B2),
				.a1(P00C2),
				.a2(P00D2),
				.a3(P01B2),
				.a4(P01C2),
				.a5(P01D2),
				.a6(P02B2),
				.a7(P02C2),
				.a8(P02D2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c020B2)
);

assign C00B2=c000B2+c010B2+c020B2;
assign A00B2=(C00B2>=0)?1:0;

ninexnine_unit ninexnine_unit_1212(
				.clk(clk),
				.rstn(rstn),
				.a0(P00C0),
				.a1(P00D0),
				.a2(P00E0),
				.a3(P01C0),
				.a4(P01D0),
				.a5(P01E0),
				.a6(P02C0),
				.a7(P02D0),
				.a8(P02E0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c000C2)
);

ninexnine_unit ninexnine_unit_1213(
				.clk(clk),
				.rstn(rstn),
				.a0(P00C1),
				.a1(P00D1),
				.a2(P00E1),
				.a3(P01C1),
				.a4(P01D1),
				.a5(P01E1),
				.a6(P02C1),
				.a7(P02D1),
				.a8(P02E1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c010C2)
);

ninexnine_unit ninexnine_unit_1214(
				.clk(clk),
				.rstn(rstn),
				.a0(P00C2),
				.a1(P00D2),
				.a2(P00E2),
				.a3(P01C2),
				.a4(P01D2),
				.a5(P01E2),
				.a6(P02C2),
				.a7(P02D2),
				.a8(P02E2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c020C2)
);

assign C00C2=c000C2+c010C2+c020C2;
assign A00C2=(C00C2>=0)?1:0;

ninexnine_unit ninexnine_unit_1215(
				.clk(clk),
				.rstn(rstn),
				.a0(P00D0),
				.a1(P00E0),
				.a2(P00F0),
				.a3(P01D0),
				.a4(P01E0),
				.a5(P01F0),
				.a6(P02D0),
				.a7(P02E0),
				.a8(P02F0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c000D2)
);

ninexnine_unit ninexnine_unit_1216(
				.clk(clk),
				.rstn(rstn),
				.a0(P00D1),
				.a1(P00E1),
				.a2(P00F1),
				.a3(P01D1),
				.a4(P01E1),
				.a5(P01F1),
				.a6(P02D1),
				.a7(P02E1),
				.a8(P02F1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c010D2)
);

ninexnine_unit ninexnine_unit_1217(
				.clk(clk),
				.rstn(rstn),
				.a0(P00D2),
				.a1(P00E2),
				.a2(P00F2),
				.a3(P01D2),
				.a4(P01E2),
				.a5(P01F2),
				.a6(P02D2),
				.a7(P02E2),
				.a8(P02F2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c020D2)
);

assign C00D2=c000D2+c010D2+c020D2;
assign A00D2=(C00D2>=0)?1:0;

ninexnine_unit ninexnine_unit_1218(
				.clk(clk),
				.rstn(rstn),
				.a0(P0100),
				.a1(P0110),
				.a2(P0120),
				.a3(P0200),
				.a4(P0210),
				.a5(P0220),
				.a6(P0300),
				.a7(P0310),
				.a8(P0320),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00102)
);

ninexnine_unit ninexnine_unit_1219(
				.clk(clk),
				.rstn(rstn),
				.a0(P0101),
				.a1(P0111),
				.a2(P0121),
				.a3(P0201),
				.a4(P0211),
				.a5(P0221),
				.a6(P0301),
				.a7(P0311),
				.a8(P0321),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01102)
);

ninexnine_unit ninexnine_unit_1220(
				.clk(clk),
				.rstn(rstn),
				.a0(P0102),
				.a1(P0112),
				.a2(P0122),
				.a3(P0202),
				.a4(P0212),
				.a5(P0222),
				.a6(P0302),
				.a7(P0312),
				.a8(P0322),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02102)
);

assign C0102=c00102+c01102+c02102;
assign A0102=(C0102>=0)?1:0;

ninexnine_unit ninexnine_unit_1221(
				.clk(clk),
				.rstn(rstn),
				.a0(P0110),
				.a1(P0120),
				.a2(P0130),
				.a3(P0210),
				.a4(P0220),
				.a5(P0230),
				.a6(P0310),
				.a7(P0320),
				.a8(P0330),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00112)
);

ninexnine_unit ninexnine_unit_1222(
				.clk(clk),
				.rstn(rstn),
				.a0(P0111),
				.a1(P0121),
				.a2(P0131),
				.a3(P0211),
				.a4(P0221),
				.a5(P0231),
				.a6(P0311),
				.a7(P0321),
				.a8(P0331),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01112)
);

ninexnine_unit ninexnine_unit_1223(
				.clk(clk),
				.rstn(rstn),
				.a0(P0112),
				.a1(P0122),
				.a2(P0132),
				.a3(P0212),
				.a4(P0222),
				.a5(P0232),
				.a6(P0312),
				.a7(P0322),
				.a8(P0332),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02112)
);

assign C0112=c00112+c01112+c02112;
assign A0112=(C0112>=0)?1:0;

ninexnine_unit ninexnine_unit_1224(
				.clk(clk),
				.rstn(rstn),
				.a0(P0120),
				.a1(P0130),
				.a2(P0140),
				.a3(P0220),
				.a4(P0230),
				.a5(P0240),
				.a6(P0320),
				.a7(P0330),
				.a8(P0340),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00122)
);

ninexnine_unit ninexnine_unit_1225(
				.clk(clk),
				.rstn(rstn),
				.a0(P0121),
				.a1(P0131),
				.a2(P0141),
				.a3(P0221),
				.a4(P0231),
				.a5(P0241),
				.a6(P0321),
				.a7(P0331),
				.a8(P0341),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01122)
);

ninexnine_unit ninexnine_unit_1226(
				.clk(clk),
				.rstn(rstn),
				.a0(P0122),
				.a1(P0132),
				.a2(P0142),
				.a3(P0222),
				.a4(P0232),
				.a5(P0242),
				.a6(P0322),
				.a7(P0332),
				.a8(P0342),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02122)
);

assign C0122=c00122+c01122+c02122;
assign A0122=(C0122>=0)?1:0;

ninexnine_unit ninexnine_unit_1227(
				.clk(clk),
				.rstn(rstn),
				.a0(P0130),
				.a1(P0140),
				.a2(P0150),
				.a3(P0230),
				.a4(P0240),
				.a5(P0250),
				.a6(P0330),
				.a7(P0340),
				.a8(P0350),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00132)
);

ninexnine_unit ninexnine_unit_1228(
				.clk(clk),
				.rstn(rstn),
				.a0(P0131),
				.a1(P0141),
				.a2(P0151),
				.a3(P0231),
				.a4(P0241),
				.a5(P0251),
				.a6(P0331),
				.a7(P0341),
				.a8(P0351),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01132)
);

ninexnine_unit ninexnine_unit_1229(
				.clk(clk),
				.rstn(rstn),
				.a0(P0132),
				.a1(P0142),
				.a2(P0152),
				.a3(P0232),
				.a4(P0242),
				.a5(P0252),
				.a6(P0332),
				.a7(P0342),
				.a8(P0352),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02132)
);

assign C0132=c00132+c01132+c02132;
assign A0132=(C0132>=0)?1:0;

ninexnine_unit ninexnine_unit_1230(
				.clk(clk),
				.rstn(rstn),
				.a0(P0140),
				.a1(P0150),
				.a2(P0160),
				.a3(P0240),
				.a4(P0250),
				.a5(P0260),
				.a6(P0340),
				.a7(P0350),
				.a8(P0360),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00142)
);

ninexnine_unit ninexnine_unit_1231(
				.clk(clk),
				.rstn(rstn),
				.a0(P0141),
				.a1(P0151),
				.a2(P0161),
				.a3(P0241),
				.a4(P0251),
				.a5(P0261),
				.a6(P0341),
				.a7(P0351),
				.a8(P0361),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01142)
);

ninexnine_unit ninexnine_unit_1232(
				.clk(clk),
				.rstn(rstn),
				.a0(P0142),
				.a1(P0152),
				.a2(P0162),
				.a3(P0242),
				.a4(P0252),
				.a5(P0262),
				.a6(P0342),
				.a7(P0352),
				.a8(P0362),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02142)
);

assign C0142=c00142+c01142+c02142;
assign A0142=(C0142>=0)?1:0;

ninexnine_unit ninexnine_unit_1233(
				.clk(clk),
				.rstn(rstn),
				.a0(P0150),
				.a1(P0160),
				.a2(P0170),
				.a3(P0250),
				.a4(P0260),
				.a5(P0270),
				.a6(P0350),
				.a7(P0360),
				.a8(P0370),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00152)
);

ninexnine_unit ninexnine_unit_1234(
				.clk(clk),
				.rstn(rstn),
				.a0(P0151),
				.a1(P0161),
				.a2(P0171),
				.a3(P0251),
				.a4(P0261),
				.a5(P0271),
				.a6(P0351),
				.a7(P0361),
				.a8(P0371),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01152)
);

ninexnine_unit ninexnine_unit_1235(
				.clk(clk),
				.rstn(rstn),
				.a0(P0152),
				.a1(P0162),
				.a2(P0172),
				.a3(P0252),
				.a4(P0262),
				.a5(P0272),
				.a6(P0352),
				.a7(P0362),
				.a8(P0372),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02152)
);

assign C0152=c00152+c01152+c02152;
assign A0152=(C0152>=0)?1:0;

ninexnine_unit ninexnine_unit_1236(
				.clk(clk),
				.rstn(rstn),
				.a0(P0160),
				.a1(P0170),
				.a2(P0180),
				.a3(P0260),
				.a4(P0270),
				.a5(P0280),
				.a6(P0360),
				.a7(P0370),
				.a8(P0380),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00162)
);

ninexnine_unit ninexnine_unit_1237(
				.clk(clk),
				.rstn(rstn),
				.a0(P0161),
				.a1(P0171),
				.a2(P0181),
				.a3(P0261),
				.a4(P0271),
				.a5(P0281),
				.a6(P0361),
				.a7(P0371),
				.a8(P0381),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01162)
);

ninexnine_unit ninexnine_unit_1238(
				.clk(clk),
				.rstn(rstn),
				.a0(P0162),
				.a1(P0172),
				.a2(P0182),
				.a3(P0262),
				.a4(P0272),
				.a5(P0282),
				.a6(P0362),
				.a7(P0372),
				.a8(P0382),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02162)
);

assign C0162=c00162+c01162+c02162;
assign A0162=(C0162>=0)?1:0;

ninexnine_unit ninexnine_unit_1239(
				.clk(clk),
				.rstn(rstn),
				.a0(P0170),
				.a1(P0180),
				.a2(P0190),
				.a3(P0270),
				.a4(P0280),
				.a5(P0290),
				.a6(P0370),
				.a7(P0380),
				.a8(P0390),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00172)
);

ninexnine_unit ninexnine_unit_1240(
				.clk(clk),
				.rstn(rstn),
				.a0(P0171),
				.a1(P0181),
				.a2(P0191),
				.a3(P0271),
				.a4(P0281),
				.a5(P0291),
				.a6(P0371),
				.a7(P0381),
				.a8(P0391),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01172)
);

ninexnine_unit ninexnine_unit_1241(
				.clk(clk),
				.rstn(rstn),
				.a0(P0172),
				.a1(P0182),
				.a2(P0192),
				.a3(P0272),
				.a4(P0282),
				.a5(P0292),
				.a6(P0372),
				.a7(P0382),
				.a8(P0392),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02172)
);

assign C0172=c00172+c01172+c02172;
assign A0172=(C0172>=0)?1:0;

ninexnine_unit ninexnine_unit_1242(
				.clk(clk),
				.rstn(rstn),
				.a0(P0180),
				.a1(P0190),
				.a2(P01A0),
				.a3(P0280),
				.a4(P0290),
				.a5(P02A0),
				.a6(P0380),
				.a7(P0390),
				.a8(P03A0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00182)
);

ninexnine_unit ninexnine_unit_1243(
				.clk(clk),
				.rstn(rstn),
				.a0(P0181),
				.a1(P0191),
				.a2(P01A1),
				.a3(P0281),
				.a4(P0291),
				.a5(P02A1),
				.a6(P0381),
				.a7(P0391),
				.a8(P03A1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01182)
);

ninexnine_unit ninexnine_unit_1244(
				.clk(clk),
				.rstn(rstn),
				.a0(P0182),
				.a1(P0192),
				.a2(P01A2),
				.a3(P0282),
				.a4(P0292),
				.a5(P02A2),
				.a6(P0382),
				.a7(P0392),
				.a8(P03A2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02182)
);

assign C0182=c00182+c01182+c02182;
assign A0182=(C0182>=0)?1:0;

ninexnine_unit ninexnine_unit_1245(
				.clk(clk),
				.rstn(rstn),
				.a0(P0190),
				.a1(P01A0),
				.a2(P01B0),
				.a3(P0290),
				.a4(P02A0),
				.a5(P02B0),
				.a6(P0390),
				.a7(P03A0),
				.a8(P03B0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00192)
);

ninexnine_unit ninexnine_unit_1246(
				.clk(clk),
				.rstn(rstn),
				.a0(P0191),
				.a1(P01A1),
				.a2(P01B1),
				.a3(P0291),
				.a4(P02A1),
				.a5(P02B1),
				.a6(P0391),
				.a7(P03A1),
				.a8(P03B1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01192)
);

ninexnine_unit ninexnine_unit_1247(
				.clk(clk),
				.rstn(rstn),
				.a0(P0192),
				.a1(P01A2),
				.a2(P01B2),
				.a3(P0292),
				.a4(P02A2),
				.a5(P02B2),
				.a6(P0392),
				.a7(P03A2),
				.a8(P03B2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02192)
);

assign C0192=c00192+c01192+c02192;
assign A0192=(C0192>=0)?1:0;

ninexnine_unit ninexnine_unit_1248(
				.clk(clk),
				.rstn(rstn),
				.a0(P01A0),
				.a1(P01B0),
				.a2(P01C0),
				.a3(P02A0),
				.a4(P02B0),
				.a5(P02C0),
				.a6(P03A0),
				.a7(P03B0),
				.a8(P03C0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c001A2)
);

ninexnine_unit ninexnine_unit_1249(
				.clk(clk),
				.rstn(rstn),
				.a0(P01A1),
				.a1(P01B1),
				.a2(P01C1),
				.a3(P02A1),
				.a4(P02B1),
				.a5(P02C1),
				.a6(P03A1),
				.a7(P03B1),
				.a8(P03C1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c011A2)
);

ninexnine_unit ninexnine_unit_1250(
				.clk(clk),
				.rstn(rstn),
				.a0(P01A2),
				.a1(P01B2),
				.a2(P01C2),
				.a3(P02A2),
				.a4(P02B2),
				.a5(P02C2),
				.a6(P03A2),
				.a7(P03B2),
				.a8(P03C2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c021A2)
);

assign C01A2=c001A2+c011A2+c021A2;
assign A01A2=(C01A2>=0)?1:0;

ninexnine_unit ninexnine_unit_1251(
				.clk(clk),
				.rstn(rstn),
				.a0(P01B0),
				.a1(P01C0),
				.a2(P01D0),
				.a3(P02B0),
				.a4(P02C0),
				.a5(P02D0),
				.a6(P03B0),
				.a7(P03C0),
				.a8(P03D0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c001B2)
);

ninexnine_unit ninexnine_unit_1252(
				.clk(clk),
				.rstn(rstn),
				.a0(P01B1),
				.a1(P01C1),
				.a2(P01D1),
				.a3(P02B1),
				.a4(P02C1),
				.a5(P02D1),
				.a6(P03B1),
				.a7(P03C1),
				.a8(P03D1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c011B2)
);

ninexnine_unit ninexnine_unit_1253(
				.clk(clk),
				.rstn(rstn),
				.a0(P01B2),
				.a1(P01C2),
				.a2(P01D2),
				.a3(P02B2),
				.a4(P02C2),
				.a5(P02D2),
				.a6(P03B2),
				.a7(P03C2),
				.a8(P03D2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c021B2)
);

assign C01B2=c001B2+c011B2+c021B2;
assign A01B2=(C01B2>=0)?1:0;

ninexnine_unit ninexnine_unit_1254(
				.clk(clk),
				.rstn(rstn),
				.a0(P01C0),
				.a1(P01D0),
				.a2(P01E0),
				.a3(P02C0),
				.a4(P02D0),
				.a5(P02E0),
				.a6(P03C0),
				.a7(P03D0),
				.a8(P03E0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c001C2)
);

ninexnine_unit ninexnine_unit_1255(
				.clk(clk),
				.rstn(rstn),
				.a0(P01C1),
				.a1(P01D1),
				.a2(P01E1),
				.a3(P02C1),
				.a4(P02D1),
				.a5(P02E1),
				.a6(P03C1),
				.a7(P03D1),
				.a8(P03E1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c011C2)
);

ninexnine_unit ninexnine_unit_1256(
				.clk(clk),
				.rstn(rstn),
				.a0(P01C2),
				.a1(P01D2),
				.a2(P01E2),
				.a3(P02C2),
				.a4(P02D2),
				.a5(P02E2),
				.a6(P03C2),
				.a7(P03D2),
				.a8(P03E2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c021C2)
);

assign C01C2=c001C2+c011C2+c021C2;
assign A01C2=(C01C2>=0)?1:0;

ninexnine_unit ninexnine_unit_1257(
				.clk(clk),
				.rstn(rstn),
				.a0(P01D0),
				.a1(P01E0),
				.a2(P01F0),
				.a3(P02D0),
				.a4(P02E0),
				.a5(P02F0),
				.a6(P03D0),
				.a7(P03E0),
				.a8(P03F0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c001D2)
);

ninexnine_unit ninexnine_unit_1258(
				.clk(clk),
				.rstn(rstn),
				.a0(P01D1),
				.a1(P01E1),
				.a2(P01F1),
				.a3(P02D1),
				.a4(P02E1),
				.a5(P02F1),
				.a6(P03D1),
				.a7(P03E1),
				.a8(P03F1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c011D2)
);

ninexnine_unit ninexnine_unit_1259(
				.clk(clk),
				.rstn(rstn),
				.a0(P01D2),
				.a1(P01E2),
				.a2(P01F2),
				.a3(P02D2),
				.a4(P02E2),
				.a5(P02F2),
				.a6(P03D2),
				.a7(P03E2),
				.a8(P03F2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c021D2)
);

assign C01D2=c001D2+c011D2+c021D2;
assign A01D2=(C01D2>=0)?1:0;

ninexnine_unit ninexnine_unit_1260(
				.clk(clk),
				.rstn(rstn),
				.a0(P0200),
				.a1(P0210),
				.a2(P0220),
				.a3(P0300),
				.a4(P0310),
				.a5(P0320),
				.a6(P0400),
				.a7(P0410),
				.a8(P0420),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00202)
);

ninexnine_unit ninexnine_unit_1261(
				.clk(clk),
				.rstn(rstn),
				.a0(P0201),
				.a1(P0211),
				.a2(P0221),
				.a3(P0301),
				.a4(P0311),
				.a5(P0321),
				.a6(P0401),
				.a7(P0411),
				.a8(P0421),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01202)
);

ninexnine_unit ninexnine_unit_1262(
				.clk(clk),
				.rstn(rstn),
				.a0(P0202),
				.a1(P0212),
				.a2(P0222),
				.a3(P0302),
				.a4(P0312),
				.a5(P0322),
				.a6(P0402),
				.a7(P0412),
				.a8(P0422),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02202)
);

assign C0202=c00202+c01202+c02202;
assign A0202=(C0202>=0)?1:0;

ninexnine_unit ninexnine_unit_1263(
				.clk(clk),
				.rstn(rstn),
				.a0(P0210),
				.a1(P0220),
				.a2(P0230),
				.a3(P0310),
				.a4(P0320),
				.a5(P0330),
				.a6(P0410),
				.a7(P0420),
				.a8(P0430),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00212)
);

ninexnine_unit ninexnine_unit_1264(
				.clk(clk),
				.rstn(rstn),
				.a0(P0211),
				.a1(P0221),
				.a2(P0231),
				.a3(P0311),
				.a4(P0321),
				.a5(P0331),
				.a6(P0411),
				.a7(P0421),
				.a8(P0431),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01212)
);

ninexnine_unit ninexnine_unit_1265(
				.clk(clk),
				.rstn(rstn),
				.a0(P0212),
				.a1(P0222),
				.a2(P0232),
				.a3(P0312),
				.a4(P0322),
				.a5(P0332),
				.a6(P0412),
				.a7(P0422),
				.a8(P0432),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02212)
);

assign C0212=c00212+c01212+c02212;
assign A0212=(C0212>=0)?1:0;

ninexnine_unit ninexnine_unit_1266(
				.clk(clk),
				.rstn(rstn),
				.a0(P0220),
				.a1(P0230),
				.a2(P0240),
				.a3(P0320),
				.a4(P0330),
				.a5(P0340),
				.a6(P0420),
				.a7(P0430),
				.a8(P0440),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00222)
);

ninexnine_unit ninexnine_unit_1267(
				.clk(clk),
				.rstn(rstn),
				.a0(P0221),
				.a1(P0231),
				.a2(P0241),
				.a3(P0321),
				.a4(P0331),
				.a5(P0341),
				.a6(P0421),
				.a7(P0431),
				.a8(P0441),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01222)
);

ninexnine_unit ninexnine_unit_1268(
				.clk(clk),
				.rstn(rstn),
				.a0(P0222),
				.a1(P0232),
				.a2(P0242),
				.a3(P0322),
				.a4(P0332),
				.a5(P0342),
				.a6(P0422),
				.a7(P0432),
				.a8(P0442),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02222)
);

assign C0222=c00222+c01222+c02222;
assign A0222=(C0222>=0)?1:0;

ninexnine_unit ninexnine_unit_1269(
				.clk(clk),
				.rstn(rstn),
				.a0(P0230),
				.a1(P0240),
				.a2(P0250),
				.a3(P0330),
				.a4(P0340),
				.a5(P0350),
				.a6(P0430),
				.a7(P0440),
				.a8(P0450),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00232)
);

ninexnine_unit ninexnine_unit_1270(
				.clk(clk),
				.rstn(rstn),
				.a0(P0231),
				.a1(P0241),
				.a2(P0251),
				.a3(P0331),
				.a4(P0341),
				.a5(P0351),
				.a6(P0431),
				.a7(P0441),
				.a8(P0451),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01232)
);

ninexnine_unit ninexnine_unit_1271(
				.clk(clk),
				.rstn(rstn),
				.a0(P0232),
				.a1(P0242),
				.a2(P0252),
				.a3(P0332),
				.a4(P0342),
				.a5(P0352),
				.a6(P0432),
				.a7(P0442),
				.a8(P0452),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02232)
);

assign C0232=c00232+c01232+c02232;
assign A0232=(C0232>=0)?1:0;

ninexnine_unit ninexnine_unit_1272(
				.clk(clk),
				.rstn(rstn),
				.a0(P0240),
				.a1(P0250),
				.a2(P0260),
				.a3(P0340),
				.a4(P0350),
				.a5(P0360),
				.a6(P0440),
				.a7(P0450),
				.a8(P0460),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00242)
);

ninexnine_unit ninexnine_unit_1273(
				.clk(clk),
				.rstn(rstn),
				.a0(P0241),
				.a1(P0251),
				.a2(P0261),
				.a3(P0341),
				.a4(P0351),
				.a5(P0361),
				.a6(P0441),
				.a7(P0451),
				.a8(P0461),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01242)
);

ninexnine_unit ninexnine_unit_1274(
				.clk(clk),
				.rstn(rstn),
				.a0(P0242),
				.a1(P0252),
				.a2(P0262),
				.a3(P0342),
				.a4(P0352),
				.a5(P0362),
				.a6(P0442),
				.a7(P0452),
				.a8(P0462),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02242)
);

assign C0242=c00242+c01242+c02242;
assign A0242=(C0242>=0)?1:0;

ninexnine_unit ninexnine_unit_1275(
				.clk(clk),
				.rstn(rstn),
				.a0(P0250),
				.a1(P0260),
				.a2(P0270),
				.a3(P0350),
				.a4(P0360),
				.a5(P0370),
				.a6(P0450),
				.a7(P0460),
				.a8(P0470),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00252)
);

ninexnine_unit ninexnine_unit_1276(
				.clk(clk),
				.rstn(rstn),
				.a0(P0251),
				.a1(P0261),
				.a2(P0271),
				.a3(P0351),
				.a4(P0361),
				.a5(P0371),
				.a6(P0451),
				.a7(P0461),
				.a8(P0471),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01252)
);

ninexnine_unit ninexnine_unit_1277(
				.clk(clk),
				.rstn(rstn),
				.a0(P0252),
				.a1(P0262),
				.a2(P0272),
				.a3(P0352),
				.a4(P0362),
				.a5(P0372),
				.a6(P0452),
				.a7(P0462),
				.a8(P0472),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02252)
);

assign C0252=c00252+c01252+c02252;
assign A0252=(C0252>=0)?1:0;

ninexnine_unit ninexnine_unit_1278(
				.clk(clk),
				.rstn(rstn),
				.a0(P0260),
				.a1(P0270),
				.a2(P0280),
				.a3(P0360),
				.a4(P0370),
				.a5(P0380),
				.a6(P0460),
				.a7(P0470),
				.a8(P0480),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00262)
);

ninexnine_unit ninexnine_unit_1279(
				.clk(clk),
				.rstn(rstn),
				.a0(P0261),
				.a1(P0271),
				.a2(P0281),
				.a3(P0361),
				.a4(P0371),
				.a5(P0381),
				.a6(P0461),
				.a7(P0471),
				.a8(P0481),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01262)
);

ninexnine_unit ninexnine_unit_1280(
				.clk(clk),
				.rstn(rstn),
				.a0(P0262),
				.a1(P0272),
				.a2(P0282),
				.a3(P0362),
				.a4(P0372),
				.a5(P0382),
				.a6(P0462),
				.a7(P0472),
				.a8(P0482),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02262)
);

assign C0262=c00262+c01262+c02262;
assign A0262=(C0262>=0)?1:0;

ninexnine_unit ninexnine_unit_1281(
				.clk(clk),
				.rstn(rstn),
				.a0(P0270),
				.a1(P0280),
				.a2(P0290),
				.a3(P0370),
				.a4(P0380),
				.a5(P0390),
				.a6(P0470),
				.a7(P0480),
				.a8(P0490),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00272)
);

ninexnine_unit ninexnine_unit_1282(
				.clk(clk),
				.rstn(rstn),
				.a0(P0271),
				.a1(P0281),
				.a2(P0291),
				.a3(P0371),
				.a4(P0381),
				.a5(P0391),
				.a6(P0471),
				.a7(P0481),
				.a8(P0491),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01272)
);

ninexnine_unit ninexnine_unit_1283(
				.clk(clk),
				.rstn(rstn),
				.a0(P0272),
				.a1(P0282),
				.a2(P0292),
				.a3(P0372),
				.a4(P0382),
				.a5(P0392),
				.a6(P0472),
				.a7(P0482),
				.a8(P0492),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02272)
);

assign C0272=c00272+c01272+c02272;
assign A0272=(C0272>=0)?1:0;

ninexnine_unit ninexnine_unit_1284(
				.clk(clk),
				.rstn(rstn),
				.a0(P0280),
				.a1(P0290),
				.a2(P02A0),
				.a3(P0380),
				.a4(P0390),
				.a5(P03A0),
				.a6(P0480),
				.a7(P0490),
				.a8(P04A0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00282)
);

ninexnine_unit ninexnine_unit_1285(
				.clk(clk),
				.rstn(rstn),
				.a0(P0281),
				.a1(P0291),
				.a2(P02A1),
				.a3(P0381),
				.a4(P0391),
				.a5(P03A1),
				.a6(P0481),
				.a7(P0491),
				.a8(P04A1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01282)
);

ninexnine_unit ninexnine_unit_1286(
				.clk(clk),
				.rstn(rstn),
				.a0(P0282),
				.a1(P0292),
				.a2(P02A2),
				.a3(P0382),
				.a4(P0392),
				.a5(P03A2),
				.a6(P0482),
				.a7(P0492),
				.a8(P04A2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02282)
);

assign C0282=c00282+c01282+c02282;
assign A0282=(C0282>=0)?1:0;

ninexnine_unit ninexnine_unit_1287(
				.clk(clk),
				.rstn(rstn),
				.a0(P0290),
				.a1(P02A0),
				.a2(P02B0),
				.a3(P0390),
				.a4(P03A0),
				.a5(P03B0),
				.a6(P0490),
				.a7(P04A0),
				.a8(P04B0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00292)
);

ninexnine_unit ninexnine_unit_1288(
				.clk(clk),
				.rstn(rstn),
				.a0(P0291),
				.a1(P02A1),
				.a2(P02B1),
				.a3(P0391),
				.a4(P03A1),
				.a5(P03B1),
				.a6(P0491),
				.a7(P04A1),
				.a8(P04B1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01292)
);

ninexnine_unit ninexnine_unit_1289(
				.clk(clk),
				.rstn(rstn),
				.a0(P0292),
				.a1(P02A2),
				.a2(P02B2),
				.a3(P0392),
				.a4(P03A2),
				.a5(P03B2),
				.a6(P0492),
				.a7(P04A2),
				.a8(P04B2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02292)
);

assign C0292=c00292+c01292+c02292;
assign A0292=(C0292>=0)?1:0;

ninexnine_unit ninexnine_unit_1290(
				.clk(clk),
				.rstn(rstn),
				.a0(P02A0),
				.a1(P02B0),
				.a2(P02C0),
				.a3(P03A0),
				.a4(P03B0),
				.a5(P03C0),
				.a6(P04A0),
				.a7(P04B0),
				.a8(P04C0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c002A2)
);

ninexnine_unit ninexnine_unit_1291(
				.clk(clk),
				.rstn(rstn),
				.a0(P02A1),
				.a1(P02B1),
				.a2(P02C1),
				.a3(P03A1),
				.a4(P03B1),
				.a5(P03C1),
				.a6(P04A1),
				.a7(P04B1),
				.a8(P04C1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c012A2)
);

ninexnine_unit ninexnine_unit_1292(
				.clk(clk),
				.rstn(rstn),
				.a0(P02A2),
				.a1(P02B2),
				.a2(P02C2),
				.a3(P03A2),
				.a4(P03B2),
				.a5(P03C2),
				.a6(P04A2),
				.a7(P04B2),
				.a8(P04C2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c022A2)
);

assign C02A2=c002A2+c012A2+c022A2;
assign A02A2=(C02A2>=0)?1:0;

ninexnine_unit ninexnine_unit_1293(
				.clk(clk),
				.rstn(rstn),
				.a0(P02B0),
				.a1(P02C0),
				.a2(P02D0),
				.a3(P03B0),
				.a4(P03C0),
				.a5(P03D0),
				.a6(P04B0),
				.a7(P04C0),
				.a8(P04D0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c002B2)
);

ninexnine_unit ninexnine_unit_1294(
				.clk(clk),
				.rstn(rstn),
				.a0(P02B1),
				.a1(P02C1),
				.a2(P02D1),
				.a3(P03B1),
				.a4(P03C1),
				.a5(P03D1),
				.a6(P04B1),
				.a7(P04C1),
				.a8(P04D1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c012B2)
);

ninexnine_unit ninexnine_unit_1295(
				.clk(clk),
				.rstn(rstn),
				.a0(P02B2),
				.a1(P02C2),
				.a2(P02D2),
				.a3(P03B2),
				.a4(P03C2),
				.a5(P03D2),
				.a6(P04B2),
				.a7(P04C2),
				.a8(P04D2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c022B2)
);

assign C02B2=c002B2+c012B2+c022B2;
assign A02B2=(C02B2>=0)?1:0;

ninexnine_unit ninexnine_unit_1296(
				.clk(clk),
				.rstn(rstn),
				.a0(P02C0),
				.a1(P02D0),
				.a2(P02E0),
				.a3(P03C0),
				.a4(P03D0),
				.a5(P03E0),
				.a6(P04C0),
				.a7(P04D0),
				.a8(P04E0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c002C2)
);

ninexnine_unit ninexnine_unit_1297(
				.clk(clk),
				.rstn(rstn),
				.a0(P02C1),
				.a1(P02D1),
				.a2(P02E1),
				.a3(P03C1),
				.a4(P03D1),
				.a5(P03E1),
				.a6(P04C1),
				.a7(P04D1),
				.a8(P04E1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c012C2)
);

ninexnine_unit ninexnine_unit_1298(
				.clk(clk),
				.rstn(rstn),
				.a0(P02C2),
				.a1(P02D2),
				.a2(P02E2),
				.a3(P03C2),
				.a4(P03D2),
				.a5(P03E2),
				.a6(P04C2),
				.a7(P04D2),
				.a8(P04E2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c022C2)
);

assign C02C2=c002C2+c012C2+c022C2;
assign A02C2=(C02C2>=0)?1:0;

ninexnine_unit ninexnine_unit_1299(
				.clk(clk),
				.rstn(rstn),
				.a0(P02D0),
				.a1(P02E0),
				.a2(P02F0),
				.a3(P03D0),
				.a4(P03E0),
				.a5(P03F0),
				.a6(P04D0),
				.a7(P04E0),
				.a8(P04F0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c002D2)
);

ninexnine_unit ninexnine_unit_1300(
				.clk(clk),
				.rstn(rstn),
				.a0(P02D1),
				.a1(P02E1),
				.a2(P02F1),
				.a3(P03D1),
				.a4(P03E1),
				.a5(P03F1),
				.a6(P04D1),
				.a7(P04E1),
				.a8(P04F1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c012D2)
);

ninexnine_unit ninexnine_unit_1301(
				.clk(clk),
				.rstn(rstn),
				.a0(P02D2),
				.a1(P02E2),
				.a2(P02F2),
				.a3(P03D2),
				.a4(P03E2),
				.a5(P03F2),
				.a6(P04D2),
				.a7(P04E2),
				.a8(P04F2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c022D2)
);

assign C02D2=c002D2+c012D2+c022D2;
assign A02D2=(C02D2>=0)?1:0;

ninexnine_unit ninexnine_unit_1302(
				.clk(clk),
				.rstn(rstn),
				.a0(P0300),
				.a1(P0310),
				.a2(P0320),
				.a3(P0400),
				.a4(P0410),
				.a5(P0420),
				.a6(P0500),
				.a7(P0510),
				.a8(P0520),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00302)
);

ninexnine_unit ninexnine_unit_1303(
				.clk(clk),
				.rstn(rstn),
				.a0(P0301),
				.a1(P0311),
				.a2(P0321),
				.a3(P0401),
				.a4(P0411),
				.a5(P0421),
				.a6(P0501),
				.a7(P0511),
				.a8(P0521),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01302)
);

ninexnine_unit ninexnine_unit_1304(
				.clk(clk),
				.rstn(rstn),
				.a0(P0302),
				.a1(P0312),
				.a2(P0322),
				.a3(P0402),
				.a4(P0412),
				.a5(P0422),
				.a6(P0502),
				.a7(P0512),
				.a8(P0522),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02302)
);

assign C0302=c00302+c01302+c02302;
assign A0302=(C0302>=0)?1:0;

ninexnine_unit ninexnine_unit_1305(
				.clk(clk),
				.rstn(rstn),
				.a0(P0310),
				.a1(P0320),
				.a2(P0330),
				.a3(P0410),
				.a4(P0420),
				.a5(P0430),
				.a6(P0510),
				.a7(P0520),
				.a8(P0530),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00312)
);

ninexnine_unit ninexnine_unit_1306(
				.clk(clk),
				.rstn(rstn),
				.a0(P0311),
				.a1(P0321),
				.a2(P0331),
				.a3(P0411),
				.a4(P0421),
				.a5(P0431),
				.a6(P0511),
				.a7(P0521),
				.a8(P0531),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01312)
);

ninexnine_unit ninexnine_unit_1307(
				.clk(clk),
				.rstn(rstn),
				.a0(P0312),
				.a1(P0322),
				.a2(P0332),
				.a3(P0412),
				.a4(P0422),
				.a5(P0432),
				.a6(P0512),
				.a7(P0522),
				.a8(P0532),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02312)
);

assign C0312=c00312+c01312+c02312;
assign A0312=(C0312>=0)?1:0;

ninexnine_unit ninexnine_unit_1308(
				.clk(clk),
				.rstn(rstn),
				.a0(P0320),
				.a1(P0330),
				.a2(P0340),
				.a3(P0420),
				.a4(P0430),
				.a5(P0440),
				.a6(P0520),
				.a7(P0530),
				.a8(P0540),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00322)
);

ninexnine_unit ninexnine_unit_1309(
				.clk(clk),
				.rstn(rstn),
				.a0(P0321),
				.a1(P0331),
				.a2(P0341),
				.a3(P0421),
				.a4(P0431),
				.a5(P0441),
				.a6(P0521),
				.a7(P0531),
				.a8(P0541),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01322)
);

ninexnine_unit ninexnine_unit_1310(
				.clk(clk),
				.rstn(rstn),
				.a0(P0322),
				.a1(P0332),
				.a2(P0342),
				.a3(P0422),
				.a4(P0432),
				.a5(P0442),
				.a6(P0522),
				.a7(P0532),
				.a8(P0542),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02322)
);

assign C0322=c00322+c01322+c02322;
assign A0322=(C0322>=0)?1:0;

ninexnine_unit ninexnine_unit_1311(
				.clk(clk),
				.rstn(rstn),
				.a0(P0330),
				.a1(P0340),
				.a2(P0350),
				.a3(P0430),
				.a4(P0440),
				.a5(P0450),
				.a6(P0530),
				.a7(P0540),
				.a8(P0550),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00332)
);

ninexnine_unit ninexnine_unit_1312(
				.clk(clk),
				.rstn(rstn),
				.a0(P0331),
				.a1(P0341),
				.a2(P0351),
				.a3(P0431),
				.a4(P0441),
				.a5(P0451),
				.a6(P0531),
				.a7(P0541),
				.a8(P0551),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01332)
);

ninexnine_unit ninexnine_unit_1313(
				.clk(clk),
				.rstn(rstn),
				.a0(P0332),
				.a1(P0342),
				.a2(P0352),
				.a3(P0432),
				.a4(P0442),
				.a5(P0452),
				.a6(P0532),
				.a7(P0542),
				.a8(P0552),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02332)
);

assign C0332=c00332+c01332+c02332;
assign A0332=(C0332>=0)?1:0;

ninexnine_unit ninexnine_unit_1314(
				.clk(clk),
				.rstn(rstn),
				.a0(P0340),
				.a1(P0350),
				.a2(P0360),
				.a3(P0440),
				.a4(P0450),
				.a5(P0460),
				.a6(P0540),
				.a7(P0550),
				.a8(P0560),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00342)
);

ninexnine_unit ninexnine_unit_1315(
				.clk(clk),
				.rstn(rstn),
				.a0(P0341),
				.a1(P0351),
				.a2(P0361),
				.a3(P0441),
				.a4(P0451),
				.a5(P0461),
				.a6(P0541),
				.a7(P0551),
				.a8(P0561),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01342)
);

ninexnine_unit ninexnine_unit_1316(
				.clk(clk),
				.rstn(rstn),
				.a0(P0342),
				.a1(P0352),
				.a2(P0362),
				.a3(P0442),
				.a4(P0452),
				.a5(P0462),
				.a6(P0542),
				.a7(P0552),
				.a8(P0562),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02342)
);

assign C0342=c00342+c01342+c02342;
assign A0342=(C0342>=0)?1:0;

ninexnine_unit ninexnine_unit_1317(
				.clk(clk),
				.rstn(rstn),
				.a0(P0350),
				.a1(P0360),
				.a2(P0370),
				.a3(P0450),
				.a4(P0460),
				.a5(P0470),
				.a6(P0550),
				.a7(P0560),
				.a8(P0570),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00352)
);

ninexnine_unit ninexnine_unit_1318(
				.clk(clk),
				.rstn(rstn),
				.a0(P0351),
				.a1(P0361),
				.a2(P0371),
				.a3(P0451),
				.a4(P0461),
				.a5(P0471),
				.a6(P0551),
				.a7(P0561),
				.a8(P0571),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01352)
);

ninexnine_unit ninexnine_unit_1319(
				.clk(clk),
				.rstn(rstn),
				.a0(P0352),
				.a1(P0362),
				.a2(P0372),
				.a3(P0452),
				.a4(P0462),
				.a5(P0472),
				.a6(P0552),
				.a7(P0562),
				.a8(P0572),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02352)
);

assign C0352=c00352+c01352+c02352;
assign A0352=(C0352>=0)?1:0;

ninexnine_unit ninexnine_unit_1320(
				.clk(clk),
				.rstn(rstn),
				.a0(P0360),
				.a1(P0370),
				.a2(P0380),
				.a3(P0460),
				.a4(P0470),
				.a5(P0480),
				.a6(P0560),
				.a7(P0570),
				.a8(P0580),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00362)
);

ninexnine_unit ninexnine_unit_1321(
				.clk(clk),
				.rstn(rstn),
				.a0(P0361),
				.a1(P0371),
				.a2(P0381),
				.a3(P0461),
				.a4(P0471),
				.a5(P0481),
				.a6(P0561),
				.a7(P0571),
				.a8(P0581),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01362)
);

ninexnine_unit ninexnine_unit_1322(
				.clk(clk),
				.rstn(rstn),
				.a0(P0362),
				.a1(P0372),
				.a2(P0382),
				.a3(P0462),
				.a4(P0472),
				.a5(P0482),
				.a6(P0562),
				.a7(P0572),
				.a8(P0582),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02362)
);

assign C0362=c00362+c01362+c02362;
assign A0362=(C0362>=0)?1:0;

ninexnine_unit ninexnine_unit_1323(
				.clk(clk),
				.rstn(rstn),
				.a0(P0370),
				.a1(P0380),
				.a2(P0390),
				.a3(P0470),
				.a4(P0480),
				.a5(P0490),
				.a6(P0570),
				.a7(P0580),
				.a8(P0590),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00372)
);

ninexnine_unit ninexnine_unit_1324(
				.clk(clk),
				.rstn(rstn),
				.a0(P0371),
				.a1(P0381),
				.a2(P0391),
				.a3(P0471),
				.a4(P0481),
				.a5(P0491),
				.a6(P0571),
				.a7(P0581),
				.a8(P0591),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01372)
);

ninexnine_unit ninexnine_unit_1325(
				.clk(clk),
				.rstn(rstn),
				.a0(P0372),
				.a1(P0382),
				.a2(P0392),
				.a3(P0472),
				.a4(P0482),
				.a5(P0492),
				.a6(P0572),
				.a7(P0582),
				.a8(P0592),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02372)
);

assign C0372=c00372+c01372+c02372;
assign A0372=(C0372>=0)?1:0;

ninexnine_unit ninexnine_unit_1326(
				.clk(clk),
				.rstn(rstn),
				.a0(P0380),
				.a1(P0390),
				.a2(P03A0),
				.a3(P0480),
				.a4(P0490),
				.a5(P04A0),
				.a6(P0580),
				.a7(P0590),
				.a8(P05A0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00382)
);

ninexnine_unit ninexnine_unit_1327(
				.clk(clk),
				.rstn(rstn),
				.a0(P0381),
				.a1(P0391),
				.a2(P03A1),
				.a3(P0481),
				.a4(P0491),
				.a5(P04A1),
				.a6(P0581),
				.a7(P0591),
				.a8(P05A1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01382)
);

ninexnine_unit ninexnine_unit_1328(
				.clk(clk),
				.rstn(rstn),
				.a0(P0382),
				.a1(P0392),
				.a2(P03A2),
				.a3(P0482),
				.a4(P0492),
				.a5(P04A2),
				.a6(P0582),
				.a7(P0592),
				.a8(P05A2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02382)
);

assign C0382=c00382+c01382+c02382;
assign A0382=(C0382>=0)?1:0;

ninexnine_unit ninexnine_unit_1329(
				.clk(clk),
				.rstn(rstn),
				.a0(P0390),
				.a1(P03A0),
				.a2(P03B0),
				.a3(P0490),
				.a4(P04A0),
				.a5(P04B0),
				.a6(P0590),
				.a7(P05A0),
				.a8(P05B0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00392)
);

ninexnine_unit ninexnine_unit_1330(
				.clk(clk),
				.rstn(rstn),
				.a0(P0391),
				.a1(P03A1),
				.a2(P03B1),
				.a3(P0491),
				.a4(P04A1),
				.a5(P04B1),
				.a6(P0591),
				.a7(P05A1),
				.a8(P05B1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01392)
);

ninexnine_unit ninexnine_unit_1331(
				.clk(clk),
				.rstn(rstn),
				.a0(P0392),
				.a1(P03A2),
				.a2(P03B2),
				.a3(P0492),
				.a4(P04A2),
				.a5(P04B2),
				.a6(P0592),
				.a7(P05A2),
				.a8(P05B2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02392)
);

assign C0392=c00392+c01392+c02392;
assign A0392=(C0392>=0)?1:0;

ninexnine_unit ninexnine_unit_1332(
				.clk(clk),
				.rstn(rstn),
				.a0(P03A0),
				.a1(P03B0),
				.a2(P03C0),
				.a3(P04A0),
				.a4(P04B0),
				.a5(P04C0),
				.a6(P05A0),
				.a7(P05B0),
				.a8(P05C0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c003A2)
);

ninexnine_unit ninexnine_unit_1333(
				.clk(clk),
				.rstn(rstn),
				.a0(P03A1),
				.a1(P03B1),
				.a2(P03C1),
				.a3(P04A1),
				.a4(P04B1),
				.a5(P04C1),
				.a6(P05A1),
				.a7(P05B1),
				.a8(P05C1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c013A2)
);

ninexnine_unit ninexnine_unit_1334(
				.clk(clk),
				.rstn(rstn),
				.a0(P03A2),
				.a1(P03B2),
				.a2(P03C2),
				.a3(P04A2),
				.a4(P04B2),
				.a5(P04C2),
				.a6(P05A2),
				.a7(P05B2),
				.a8(P05C2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c023A2)
);

assign C03A2=c003A2+c013A2+c023A2;
assign A03A2=(C03A2>=0)?1:0;

ninexnine_unit ninexnine_unit_1335(
				.clk(clk),
				.rstn(rstn),
				.a0(P03B0),
				.a1(P03C0),
				.a2(P03D0),
				.a3(P04B0),
				.a4(P04C0),
				.a5(P04D0),
				.a6(P05B0),
				.a7(P05C0),
				.a8(P05D0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c003B2)
);

ninexnine_unit ninexnine_unit_1336(
				.clk(clk),
				.rstn(rstn),
				.a0(P03B1),
				.a1(P03C1),
				.a2(P03D1),
				.a3(P04B1),
				.a4(P04C1),
				.a5(P04D1),
				.a6(P05B1),
				.a7(P05C1),
				.a8(P05D1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c013B2)
);

ninexnine_unit ninexnine_unit_1337(
				.clk(clk),
				.rstn(rstn),
				.a0(P03B2),
				.a1(P03C2),
				.a2(P03D2),
				.a3(P04B2),
				.a4(P04C2),
				.a5(P04D2),
				.a6(P05B2),
				.a7(P05C2),
				.a8(P05D2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c023B2)
);

assign C03B2=c003B2+c013B2+c023B2;
assign A03B2=(C03B2>=0)?1:0;

ninexnine_unit ninexnine_unit_1338(
				.clk(clk),
				.rstn(rstn),
				.a0(P03C0),
				.a1(P03D0),
				.a2(P03E0),
				.a3(P04C0),
				.a4(P04D0),
				.a5(P04E0),
				.a6(P05C0),
				.a7(P05D0),
				.a8(P05E0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c003C2)
);

ninexnine_unit ninexnine_unit_1339(
				.clk(clk),
				.rstn(rstn),
				.a0(P03C1),
				.a1(P03D1),
				.a2(P03E1),
				.a3(P04C1),
				.a4(P04D1),
				.a5(P04E1),
				.a6(P05C1),
				.a7(P05D1),
				.a8(P05E1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c013C2)
);

ninexnine_unit ninexnine_unit_1340(
				.clk(clk),
				.rstn(rstn),
				.a0(P03C2),
				.a1(P03D2),
				.a2(P03E2),
				.a3(P04C2),
				.a4(P04D2),
				.a5(P04E2),
				.a6(P05C2),
				.a7(P05D2),
				.a8(P05E2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c023C2)
);

assign C03C2=c003C2+c013C2+c023C2;
assign A03C2=(C03C2>=0)?1:0;

ninexnine_unit ninexnine_unit_1341(
				.clk(clk),
				.rstn(rstn),
				.a0(P03D0),
				.a1(P03E0),
				.a2(P03F0),
				.a3(P04D0),
				.a4(P04E0),
				.a5(P04F0),
				.a6(P05D0),
				.a7(P05E0),
				.a8(P05F0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c003D2)
);

ninexnine_unit ninexnine_unit_1342(
				.clk(clk),
				.rstn(rstn),
				.a0(P03D1),
				.a1(P03E1),
				.a2(P03F1),
				.a3(P04D1),
				.a4(P04E1),
				.a5(P04F1),
				.a6(P05D1),
				.a7(P05E1),
				.a8(P05F1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c013D2)
);

ninexnine_unit ninexnine_unit_1343(
				.clk(clk),
				.rstn(rstn),
				.a0(P03D2),
				.a1(P03E2),
				.a2(P03F2),
				.a3(P04D2),
				.a4(P04E2),
				.a5(P04F2),
				.a6(P05D2),
				.a7(P05E2),
				.a8(P05F2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c023D2)
);

assign C03D2=c003D2+c013D2+c023D2;
assign A03D2=(C03D2>=0)?1:0;

ninexnine_unit ninexnine_unit_1344(
				.clk(clk),
				.rstn(rstn),
				.a0(P0400),
				.a1(P0410),
				.a2(P0420),
				.a3(P0500),
				.a4(P0510),
				.a5(P0520),
				.a6(P0600),
				.a7(P0610),
				.a8(P0620),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00402)
);

ninexnine_unit ninexnine_unit_1345(
				.clk(clk),
				.rstn(rstn),
				.a0(P0401),
				.a1(P0411),
				.a2(P0421),
				.a3(P0501),
				.a4(P0511),
				.a5(P0521),
				.a6(P0601),
				.a7(P0611),
				.a8(P0621),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01402)
);

ninexnine_unit ninexnine_unit_1346(
				.clk(clk),
				.rstn(rstn),
				.a0(P0402),
				.a1(P0412),
				.a2(P0422),
				.a3(P0502),
				.a4(P0512),
				.a5(P0522),
				.a6(P0602),
				.a7(P0612),
				.a8(P0622),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02402)
);

assign C0402=c00402+c01402+c02402;
assign A0402=(C0402>=0)?1:0;

ninexnine_unit ninexnine_unit_1347(
				.clk(clk),
				.rstn(rstn),
				.a0(P0410),
				.a1(P0420),
				.a2(P0430),
				.a3(P0510),
				.a4(P0520),
				.a5(P0530),
				.a6(P0610),
				.a7(P0620),
				.a8(P0630),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00412)
);

ninexnine_unit ninexnine_unit_1348(
				.clk(clk),
				.rstn(rstn),
				.a0(P0411),
				.a1(P0421),
				.a2(P0431),
				.a3(P0511),
				.a4(P0521),
				.a5(P0531),
				.a6(P0611),
				.a7(P0621),
				.a8(P0631),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01412)
);

ninexnine_unit ninexnine_unit_1349(
				.clk(clk),
				.rstn(rstn),
				.a0(P0412),
				.a1(P0422),
				.a2(P0432),
				.a3(P0512),
				.a4(P0522),
				.a5(P0532),
				.a6(P0612),
				.a7(P0622),
				.a8(P0632),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02412)
);

assign C0412=c00412+c01412+c02412;
assign A0412=(C0412>=0)?1:0;

ninexnine_unit ninexnine_unit_1350(
				.clk(clk),
				.rstn(rstn),
				.a0(P0420),
				.a1(P0430),
				.a2(P0440),
				.a3(P0520),
				.a4(P0530),
				.a5(P0540),
				.a6(P0620),
				.a7(P0630),
				.a8(P0640),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00422)
);

ninexnine_unit ninexnine_unit_1351(
				.clk(clk),
				.rstn(rstn),
				.a0(P0421),
				.a1(P0431),
				.a2(P0441),
				.a3(P0521),
				.a4(P0531),
				.a5(P0541),
				.a6(P0621),
				.a7(P0631),
				.a8(P0641),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01422)
);

ninexnine_unit ninexnine_unit_1352(
				.clk(clk),
				.rstn(rstn),
				.a0(P0422),
				.a1(P0432),
				.a2(P0442),
				.a3(P0522),
				.a4(P0532),
				.a5(P0542),
				.a6(P0622),
				.a7(P0632),
				.a8(P0642),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02422)
);

assign C0422=c00422+c01422+c02422;
assign A0422=(C0422>=0)?1:0;

ninexnine_unit ninexnine_unit_1353(
				.clk(clk),
				.rstn(rstn),
				.a0(P0430),
				.a1(P0440),
				.a2(P0450),
				.a3(P0530),
				.a4(P0540),
				.a5(P0550),
				.a6(P0630),
				.a7(P0640),
				.a8(P0650),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00432)
);

ninexnine_unit ninexnine_unit_1354(
				.clk(clk),
				.rstn(rstn),
				.a0(P0431),
				.a1(P0441),
				.a2(P0451),
				.a3(P0531),
				.a4(P0541),
				.a5(P0551),
				.a6(P0631),
				.a7(P0641),
				.a8(P0651),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01432)
);

ninexnine_unit ninexnine_unit_1355(
				.clk(clk),
				.rstn(rstn),
				.a0(P0432),
				.a1(P0442),
				.a2(P0452),
				.a3(P0532),
				.a4(P0542),
				.a5(P0552),
				.a6(P0632),
				.a7(P0642),
				.a8(P0652),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02432)
);

assign C0432=c00432+c01432+c02432;
assign A0432=(C0432>=0)?1:0;

ninexnine_unit ninexnine_unit_1356(
				.clk(clk),
				.rstn(rstn),
				.a0(P0440),
				.a1(P0450),
				.a2(P0460),
				.a3(P0540),
				.a4(P0550),
				.a5(P0560),
				.a6(P0640),
				.a7(P0650),
				.a8(P0660),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00442)
);

ninexnine_unit ninexnine_unit_1357(
				.clk(clk),
				.rstn(rstn),
				.a0(P0441),
				.a1(P0451),
				.a2(P0461),
				.a3(P0541),
				.a4(P0551),
				.a5(P0561),
				.a6(P0641),
				.a7(P0651),
				.a8(P0661),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01442)
);

ninexnine_unit ninexnine_unit_1358(
				.clk(clk),
				.rstn(rstn),
				.a0(P0442),
				.a1(P0452),
				.a2(P0462),
				.a3(P0542),
				.a4(P0552),
				.a5(P0562),
				.a6(P0642),
				.a7(P0652),
				.a8(P0662),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02442)
);

assign C0442=c00442+c01442+c02442;
assign A0442=(C0442>=0)?1:0;

ninexnine_unit ninexnine_unit_1359(
				.clk(clk),
				.rstn(rstn),
				.a0(P0450),
				.a1(P0460),
				.a2(P0470),
				.a3(P0550),
				.a4(P0560),
				.a5(P0570),
				.a6(P0650),
				.a7(P0660),
				.a8(P0670),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00452)
);

ninexnine_unit ninexnine_unit_1360(
				.clk(clk),
				.rstn(rstn),
				.a0(P0451),
				.a1(P0461),
				.a2(P0471),
				.a3(P0551),
				.a4(P0561),
				.a5(P0571),
				.a6(P0651),
				.a7(P0661),
				.a8(P0671),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01452)
);

ninexnine_unit ninexnine_unit_1361(
				.clk(clk),
				.rstn(rstn),
				.a0(P0452),
				.a1(P0462),
				.a2(P0472),
				.a3(P0552),
				.a4(P0562),
				.a5(P0572),
				.a6(P0652),
				.a7(P0662),
				.a8(P0672),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02452)
);

assign C0452=c00452+c01452+c02452;
assign A0452=(C0452>=0)?1:0;

ninexnine_unit ninexnine_unit_1362(
				.clk(clk),
				.rstn(rstn),
				.a0(P0460),
				.a1(P0470),
				.a2(P0480),
				.a3(P0560),
				.a4(P0570),
				.a5(P0580),
				.a6(P0660),
				.a7(P0670),
				.a8(P0680),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00462)
);

ninexnine_unit ninexnine_unit_1363(
				.clk(clk),
				.rstn(rstn),
				.a0(P0461),
				.a1(P0471),
				.a2(P0481),
				.a3(P0561),
				.a4(P0571),
				.a5(P0581),
				.a6(P0661),
				.a7(P0671),
				.a8(P0681),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01462)
);

ninexnine_unit ninexnine_unit_1364(
				.clk(clk),
				.rstn(rstn),
				.a0(P0462),
				.a1(P0472),
				.a2(P0482),
				.a3(P0562),
				.a4(P0572),
				.a5(P0582),
				.a6(P0662),
				.a7(P0672),
				.a8(P0682),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02462)
);

assign C0462=c00462+c01462+c02462;
assign A0462=(C0462>=0)?1:0;

ninexnine_unit ninexnine_unit_1365(
				.clk(clk),
				.rstn(rstn),
				.a0(P0470),
				.a1(P0480),
				.a2(P0490),
				.a3(P0570),
				.a4(P0580),
				.a5(P0590),
				.a6(P0670),
				.a7(P0680),
				.a8(P0690),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00472)
);

ninexnine_unit ninexnine_unit_1366(
				.clk(clk),
				.rstn(rstn),
				.a0(P0471),
				.a1(P0481),
				.a2(P0491),
				.a3(P0571),
				.a4(P0581),
				.a5(P0591),
				.a6(P0671),
				.a7(P0681),
				.a8(P0691),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01472)
);

ninexnine_unit ninexnine_unit_1367(
				.clk(clk),
				.rstn(rstn),
				.a0(P0472),
				.a1(P0482),
				.a2(P0492),
				.a3(P0572),
				.a4(P0582),
				.a5(P0592),
				.a6(P0672),
				.a7(P0682),
				.a8(P0692),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02472)
);

assign C0472=c00472+c01472+c02472;
assign A0472=(C0472>=0)?1:0;

ninexnine_unit ninexnine_unit_1368(
				.clk(clk),
				.rstn(rstn),
				.a0(P0480),
				.a1(P0490),
				.a2(P04A0),
				.a3(P0580),
				.a4(P0590),
				.a5(P05A0),
				.a6(P0680),
				.a7(P0690),
				.a8(P06A0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00482)
);

ninexnine_unit ninexnine_unit_1369(
				.clk(clk),
				.rstn(rstn),
				.a0(P0481),
				.a1(P0491),
				.a2(P04A1),
				.a3(P0581),
				.a4(P0591),
				.a5(P05A1),
				.a6(P0681),
				.a7(P0691),
				.a8(P06A1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01482)
);

ninexnine_unit ninexnine_unit_1370(
				.clk(clk),
				.rstn(rstn),
				.a0(P0482),
				.a1(P0492),
				.a2(P04A2),
				.a3(P0582),
				.a4(P0592),
				.a5(P05A2),
				.a6(P0682),
				.a7(P0692),
				.a8(P06A2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02482)
);

assign C0482=c00482+c01482+c02482;
assign A0482=(C0482>=0)?1:0;

ninexnine_unit ninexnine_unit_1371(
				.clk(clk),
				.rstn(rstn),
				.a0(P0490),
				.a1(P04A0),
				.a2(P04B0),
				.a3(P0590),
				.a4(P05A0),
				.a5(P05B0),
				.a6(P0690),
				.a7(P06A0),
				.a8(P06B0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00492)
);

ninexnine_unit ninexnine_unit_1372(
				.clk(clk),
				.rstn(rstn),
				.a0(P0491),
				.a1(P04A1),
				.a2(P04B1),
				.a3(P0591),
				.a4(P05A1),
				.a5(P05B1),
				.a6(P0691),
				.a7(P06A1),
				.a8(P06B1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01492)
);

ninexnine_unit ninexnine_unit_1373(
				.clk(clk),
				.rstn(rstn),
				.a0(P0492),
				.a1(P04A2),
				.a2(P04B2),
				.a3(P0592),
				.a4(P05A2),
				.a5(P05B2),
				.a6(P0692),
				.a7(P06A2),
				.a8(P06B2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02492)
);

assign C0492=c00492+c01492+c02492;
assign A0492=(C0492>=0)?1:0;

ninexnine_unit ninexnine_unit_1374(
				.clk(clk),
				.rstn(rstn),
				.a0(P04A0),
				.a1(P04B0),
				.a2(P04C0),
				.a3(P05A0),
				.a4(P05B0),
				.a5(P05C0),
				.a6(P06A0),
				.a7(P06B0),
				.a8(P06C0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c004A2)
);

ninexnine_unit ninexnine_unit_1375(
				.clk(clk),
				.rstn(rstn),
				.a0(P04A1),
				.a1(P04B1),
				.a2(P04C1),
				.a3(P05A1),
				.a4(P05B1),
				.a5(P05C1),
				.a6(P06A1),
				.a7(P06B1),
				.a8(P06C1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c014A2)
);

ninexnine_unit ninexnine_unit_1376(
				.clk(clk),
				.rstn(rstn),
				.a0(P04A2),
				.a1(P04B2),
				.a2(P04C2),
				.a3(P05A2),
				.a4(P05B2),
				.a5(P05C2),
				.a6(P06A2),
				.a7(P06B2),
				.a8(P06C2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c024A2)
);

assign C04A2=c004A2+c014A2+c024A2;
assign A04A2=(C04A2>=0)?1:0;

ninexnine_unit ninexnine_unit_1377(
				.clk(clk),
				.rstn(rstn),
				.a0(P04B0),
				.a1(P04C0),
				.a2(P04D0),
				.a3(P05B0),
				.a4(P05C0),
				.a5(P05D0),
				.a6(P06B0),
				.a7(P06C0),
				.a8(P06D0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c004B2)
);

ninexnine_unit ninexnine_unit_1378(
				.clk(clk),
				.rstn(rstn),
				.a0(P04B1),
				.a1(P04C1),
				.a2(P04D1),
				.a3(P05B1),
				.a4(P05C1),
				.a5(P05D1),
				.a6(P06B1),
				.a7(P06C1),
				.a8(P06D1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c014B2)
);

ninexnine_unit ninexnine_unit_1379(
				.clk(clk),
				.rstn(rstn),
				.a0(P04B2),
				.a1(P04C2),
				.a2(P04D2),
				.a3(P05B2),
				.a4(P05C2),
				.a5(P05D2),
				.a6(P06B2),
				.a7(P06C2),
				.a8(P06D2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c024B2)
);

assign C04B2=c004B2+c014B2+c024B2;
assign A04B2=(C04B2>=0)?1:0;

ninexnine_unit ninexnine_unit_1380(
				.clk(clk),
				.rstn(rstn),
				.a0(P04C0),
				.a1(P04D0),
				.a2(P04E0),
				.a3(P05C0),
				.a4(P05D0),
				.a5(P05E0),
				.a6(P06C0),
				.a7(P06D0),
				.a8(P06E0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c004C2)
);

ninexnine_unit ninexnine_unit_1381(
				.clk(clk),
				.rstn(rstn),
				.a0(P04C1),
				.a1(P04D1),
				.a2(P04E1),
				.a3(P05C1),
				.a4(P05D1),
				.a5(P05E1),
				.a6(P06C1),
				.a7(P06D1),
				.a8(P06E1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c014C2)
);

ninexnine_unit ninexnine_unit_1382(
				.clk(clk),
				.rstn(rstn),
				.a0(P04C2),
				.a1(P04D2),
				.a2(P04E2),
				.a3(P05C2),
				.a4(P05D2),
				.a5(P05E2),
				.a6(P06C2),
				.a7(P06D2),
				.a8(P06E2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c024C2)
);

assign C04C2=c004C2+c014C2+c024C2;
assign A04C2=(C04C2>=0)?1:0;

ninexnine_unit ninexnine_unit_1383(
				.clk(clk),
				.rstn(rstn),
				.a0(P04D0),
				.a1(P04E0),
				.a2(P04F0),
				.a3(P05D0),
				.a4(P05E0),
				.a5(P05F0),
				.a6(P06D0),
				.a7(P06E0),
				.a8(P06F0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c004D2)
);

ninexnine_unit ninexnine_unit_1384(
				.clk(clk),
				.rstn(rstn),
				.a0(P04D1),
				.a1(P04E1),
				.a2(P04F1),
				.a3(P05D1),
				.a4(P05E1),
				.a5(P05F1),
				.a6(P06D1),
				.a7(P06E1),
				.a8(P06F1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c014D2)
);

ninexnine_unit ninexnine_unit_1385(
				.clk(clk),
				.rstn(rstn),
				.a0(P04D2),
				.a1(P04E2),
				.a2(P04F2),
				.a3(P05D2),
				.a4(P05E2),
				.a5(P05F2),
				.a6(P06D2),
				.a7(P06E2),
				.a8(P06F2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c024D2)
);

assign C04D2=c004D2+c014D2+c024D2;
assign A04D2=(C04D2>=0)?1:0;

ninexnine_unit ninexnine_unit_1386(
				.clk(clk),
				.rstn(rstn),
				.a0(P0500),
				.a1(P0510),
				.a2(P0520),
				.a3(P0600),
				.a4(P0610),
				.a5(P0620),
				.a6(P0700),
				.a7(P0710),
				.a8(P0720),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00502)
);

ninexnine_unit ninexnine_unit_1387(
				.clk(clk),
				.rstn(rstn),
				.a0(P0501),
				.a1(P0511),
				.a2(P0521),
				.a3(P0601),
				.a4(P0611),
				.a5(P0621),
				.a6(P0701),
				.a7(P0711),
				.a8(P0721),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01502)
);

ninexnine_unit ninexnine_unit_1388(
				.clk(clk),
				.rstn(rstn),
				.a0(P0502),
				.a1(P0512),
				.a2(P0522),
				.a3(P0602),
				.a4(P0612),
				.a5(P0622),
				.a6(P0702),
				.a7(P0712),
				.a8(P0722),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02502)
);

assign C0502=c00502+c01502+c02502;
assign A0502=(C0502>=0)?1:0;

ninexnine_unit ninexnine_unit_1389(
				.clk(clk),
				.rstn(rstn),
				.a0(P0510),
				.a1(P0520),
				.a2(P0530),
				.a3(P0610),
				.a4(P0620),
				.a5(P0630),
				.a6(P0710),
				.a7(P0720),
				.a8(P0730),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00512)
);

ninexnine_unit ninexnine_unit_1390(
				.clk(clk),
				.rstn(rstn),
				.a0(P0511),
				.a1(P0521),
				.a2(P0531),
				.a3(P0611),
				.a4(P0621),
				.a5(P0631),
				.a6(P0711),
				.a7(P0721),
				.a8(P0731),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01512)
);

ninexnine_unit ninexnine_unit_1391(
				.clk(clk),
				.rstn(rstn),
				.a0(P0512),
				.a1(P0522),
				.a2(P0532),
				.a3(P0612),
				.a4(P0622),
				.a5(P0632),
				.a6(P0712),
				.a7(P0722),
				.a8(P0732),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02512)
);

assign C0512=c00512+c01512+c02512;
assign A0512=(C0512>=0)?1:0;

ninexnine_unit ninexnine_unit_1392(
				.clk(clk),
				.rstn(rstn),
				.a0(P0520),
				.a1(P0530),
				.a2(P0540),
				.a3(P0620),
				.a4(P0630),
				.a5(P0640),
				.a6(P0720),
				.a7(P0730),
				.a8(P0740),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00522)
);

ninexnine_unit ninexnine_unit_1393(
				.clk(clk),
				.rstn(rstn),
				.a0(P0521),
				.a1(P0531),
				.a2(P0541),
				.a3(P0621),
				.a4(P0631),
				.a5(P0641),
				.a6(P0721),
				.a7(P0731),
				.a8(P0741),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01522)
);

ninexnine_unit ninexnine_unit_1394(
				.clk(clk),
				.rstn(rstn),
				.a0(P0522),
				.a1(P0532),
				.a2(P0542),
				.a3(P0622),
				.a4(P0632),
				.a5(P0642),
				.a6(P0722),
				.a7(P0732),
				.a8(P0742),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02522)
);

assign C0522=c00522+c01522+c02522;
assign A0522=(C0522>=0)?1:0;

ninexnine_unit ninexnine_unit_1395(
				.clk(clk),
				.rstn(rstn),
				.a0(P0530),
				.a1(P0540),
				.a2(P0550),
				.a3(P0630),
				.a4(P0640),
				.a5(P0650),
				.a6(P0730),
				.a7(P0740),
				.a8(P0750),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00532)
);

ninexnine_unit ninexnine_unit_1396(
				.clk(clk),
				.rstn(rstn),
				.a0(P0531),
				.a1(P0541),
				.a2(P0551),
				.a3(P0631),
				.a4(P0641),
				.a5(P0651),
				.a6(P0731),
				.a7(P0741),
				.a8(P0751),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01532)
);

ninexnine_unit ninexnine_unit_1397(
				.clk(clk),
				.rstn(rstn),
				.a0(P0532),
				.a1(P0542),
				.a2(P0552),
				.a3(P0632),
				.a4(P0642),
				.a5(P0652),
				.a6(P0732),
				.a7(P0742),
				.a8(P0752),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02532)
);

assign C0532=c00532+c01532+c02532;
assign A0532=(C0532>=0)?1:0;

ninexnine_unit ninexnine_unit_1398(
				.clk(clk),
				.rstn(rstn),
				.a0(P0540),
				.a1(P0550),
				.a2(P0560),
				.a3(P0640),
				.a4(P0650),
				.a5(P0660),
				.a6(P0740),
				.a7(P0750),
				.a8(P0760),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00542)
);

ninexnine_unit ninexnine_unit_1399(
				.clk(clk),
				.rstn(rstn),
				.a0(P0541),
				.a1(P0551),
				.a2(P0561),
				.a3(P0641),
				.a4(P0651),
				.a5(P0661),
				.a6(P0741),
				.a7(P0751),
				.a8(P0761),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01542)
);

ninexnine_unit ninexnine_unit_1400(
				.clk(clk),
				.rstn(rstn),
				.a0(P0542),
				.a1(P0552),
				.a2(P0562),
				.a3(P0642),
				.a4(P0652),
				.a5(P0662),
				.a6(P0742),
				.a7(P0752),
				.a8(P0762),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02542)
);

assign C0542=c00542+c01542+c02542;
assign A0542=(C0542>=0)?1:0;

ninexnine_unit ninexnine_unit_1401(
				.clk(clk),
				.rstn(rstn),
				.a0(P0550),
				.a1(P0560),
				.a2(P0570),
				.a3(P0650),
				.a4(P0660),
				.a5(P0670),
				.a6(P0750),
				.a7(P0760),
				.a8(P0770),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00552)
);

ninexnine_unit ninexnine_unit_1402(
				.clk(clk),
				.rstn(rstn),
				.a0(P0551),
				.a1(P0561),
				.a2(P0571),
				.a3(P0651),
				.a4(P0661),
				.a5(P0671),
				.a6(P0751),
				.a7(P0761),
				.a8(P0771),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01552)
);

ninexnine_unit ninexnine_unit_1403(
				.clk(clk),
				.rstn(rstn),
				.a0(P0552),
				.a1(P0562),
				.a2(P0572),
				.a3(P0652),
				.a4(P0662),
				.a5(P0672),
				.a6(P0752),
				.a7(P0762),
				.a8(P0772),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02552)
);

assign C0552=c00552+c01552+c02552;
assign A0552=(C0552>=0)?1:0;

ninexnine_unit ninexnine_unit_1404(
				.clk(clk),
				.rstn(rstn),
				.a0(P0560),
				.a1(P0570),
				.a2(P0580),
				.a3(P0660),
				.a4(P0670),
				.a5(P0680),
				.a6(P0760),
				.a7(P0770),
				.a8(P0780),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00562)
);

ninexnine_unit ninexnine_unit_1405(
				.clk(clk),
				.rstn(rstn),
				.a0(P0561),
				.a1(P0571),
				.a2(P0581),
				.a3(P0661),
				.a4(P0671),
				.a5(P0681),
				.a6(P0761),
				.a7(P0771),
				.a8(P0781),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01562)
);

ninexnine_unit ninexnine_unit_1406(
				.clk(clk),
				.rstn(rstn),
				.a0(P0562),
				.a1(P0572),
				.a2(P0582),
				.a3(P0662),
				.a4(P0672),
				.a5(P0682),
				.a6(P0762),
				.a7(P0772),
				.a8(P0782),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02562)
);

assign C0562=c00562+c01562+c02562;
assign A0562=(C0562>=0)?1:0;

ninexnine_unit ninexnine_unit_1407(
				.clk(clk),
				.rstn(rstn),
				.a0(P0570),
				.a1(P0580),
				.a2(P0590),
				.a3(P0670),
				.a4(P0680),
				.a5(P0690),
				.a6(P0770),
				.a7(P0780),
				.a8(P0790),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00572)
);

ninexnine_unit ninexnine_unit_1408(
				.clk(clk),
				.rstn(rstn),
				.a0(P0571),
				.a1(P0581),
				.a2(P0591),
				.a3(P0671),
				.a4(P0681),
				.a5(P0691),
				.a6(P0771),
				.a7(P0781),
				.a8(P0791),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01572)
);

ninexnine_unit ninexnine_unit_1409(
				.clk(clk),
				.rstn(rstn),
				.a0(P0572),
				.a1(P0582),
				.a2(P0592),
				.a3(P0672),
				.a4(P0682),
				.a5(P0692),
				.a6(P0772),
				.a7(P0782),
				.a8(P0792),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02572)
);

assign C0572=c00572+c01572+c02572;
assign A0572=(C0572>=0)?1:0;

ninexnine_unit ninexnine_unit_1410(
				.clk(clk),
				.rstn(rstn),
				.a0(P0580),
				.a1(P0590),
				.a2(P05A0),
				.a3(P0680),
				.a4(P0690),
				.a5(P06A0),
				.a6(P0780),
				.a7(P0790),
				.a8(P07A0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00582)
);

ninexnine_unit ninexnine_unit_1411(
				.clk(clk),
				.rstn(rstn),
				.a0(P0581),
				.a1(P0591),
				.a2(P05A1),
				.a3(P0681),
				.a4(P0691),
				.a5(P06A1),
				.a6(P0781),
				.a7(P0791),
				.a8(P07A1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01582)
);

ninexnine_unit ninexnine_unit_1412(
				.clk(clk),
				.rstn(rstn),
				.a0(P0582),
				.a1(P0592),
				.a2(P05A2),
				.a3(P0682),
				.a4(P0692),
				.a5(P06A2),
				.a6(P0782),
				.a7(P0792),
				.a8(P07A2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02582)
);

assign C0582=c00582+c01582+c02582;
assign A0582=(C0582>=0)?1:0;

ninexnine_unit ninexnine_unit_1413(
				.clk(clk),
				.rstn(rstn),
				.a0(P0590),
				.a1(P05A0),
				.a2(P05B0),
				.a3(P0690),
				.a4(P06A0),
				.a5(P06B0),
				.a6(P0790),
				.a7(P07A0),
				.a8(P07B0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00592)
);

ninexnine_unit ninexnine_unit_1414(
				.clk(clk),
				.rstn(rstn),
				.a0(P0591),
				.a1(P05A1),
				.a2(P05B1),
				.a3(P0691),
				.a4(P06A1),
				.a5(P06B1),
				.a6(P0791),
				.a7(P07A1),
				.a8(P07B1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01592)
);

ninexnine_unit ninexnine_unit_1415(
				.clk(clk),
				.rstn(rstn),
				.a0(P0592),
				.a1(P05A2),
				.a2(P05B2),
				.a3(P0692),
				.a4(P06A2),
				.a5(P06B2),
				.a6(P0792),
				.a7(P07A2),
				.a8(P07B2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02592)
);

assign C0592=c00592+c01592+c02592;
assign A0592=(C0592>=0)?1:0;

ninexnine_unit ninexnine_unit_1416(
				.clk(clk),
				.rstn(rstn),
				.a0(P05A0),
				.a1(P05B0),
				.a2(P05C0),
				.a3(P06A0),
				.a4(P06B0),
				.a5(P06C0),
				.a6(P07A0),
				.a7(P07B0),
				.a8(P07C0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c005A2)
);

ninexnine_unit ninexnine_unit_1417(
				.clk(clk),
				.rstn(rstn),
				.a0(P05A1),
				.a1(P05B1),
				.a2(P05C1),
				.a3(P06A1),
				.a4(P06B1),
				.a5(P06C1),
				.a6(P07A1),
				.a7(P07B1),
				.a8(P07C1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c015A2)
);

ninexnine_unit ninexnine_unit_1418(
				.clk(clk),
				.rstn(rstn),
				.a0(P05A2),
				.a1(P05B2),
				.a2(P05C2),
				.a3(P06A2),
				.a4(P06B2),
				.a5(P06C2),
				.a6(P07A2),
				.a7(P07B2),
				.a8(P07C2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c025A2)
);

assign C05A2=c005A2+c015A2+c025A2;
assign A05A2=(C05A2>=0)?1:0;

ninexnine_unit ninexnine_unit_1419(
				.clk(clk),
				.rstn(rstn),
				.a0(P05B0),
				.a1(P05C0),
				.a2(P05D0),
				.a3(P06B0),
				.a4(P06C0),
				.a5(P06D0),
				.a6(P07B0),
				.a7(P07C0),
				.a8(P07D0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c005B2)
);

ninexnine_unit ninexnine_unit_1420(
				.clk(clk),
				.rstn(rstn),
				.a0(P05B1),
				.a1(P05C1),
				.a2(P05D1),
				.a3(P06B1),
				.a4(P06C1),
				.a5(P06D1),
				.a6(P07B1),
				.a7(P07C1),
				.a8(P07D1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c015B2)
);

ninexnine_unit ninexnine_unit_1421(
				.clk(clk),
				.rstn(rstn),
				.a0(P05B2),
				.a1(P05C2),
				.a2(P05D2),
				.a3(P06B2),
				.a4(P06C2),
				.a5(P06D2),
				.a6(P07B2),
				.a7(P07C2),
				.a8(P07D2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c025B2)
);

assign C05B2=c005B2+c015B2+c025B2;
assign A05B2=(C05B2>=0)?1:0;

ninexnine_unit ninexnine_unit_1422(
				.clk(clk),
				.rstn(rstn),
				.a0(P05C0),
				.a1(P05D0),
				.a2(P05E0),
				.a3(P06C0),
				.a4(P06D0),
				.a5(P06E0),
				.a6(P07C0),
				.a7(P07D0),
				.a8(P07E0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c005C2)
);

ninexnine_unit ninexnine_unit_1423(
				.clk(clk),
				.rstn(rstn),
				.a0(P05C1),
				.a1(P05D1),
				.a2(P05E1),
				.a3(P06C1),
				.a4(P06D1),
				.a5(P06E1),
				.a6(P07C1),
				.a7(P07D1),
				.a8(P07E1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c015C2)
);

ninexnine_unit ninexnine_unit_1424(
				.clk(clk),
				.rstn(rstn),
				.a0(P05C2),
				.a1(P05D2),
				.a2(P05E2),
				.a3(P06C2),
				.a4(P06D2),
				.a5(P06E2),
				.a6(P07C2),
				.a7(P07D2),
				.a8(P07E2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c025C2)
);

assign C05C2=c005C2+c015C2+c025C2;
assign A05C2=(C05C2>=0)?1:0;

ninexnine_unit ninexnine_unit_1425(
				.clk(clk),
				.rstn(rstn),
				.a0(P05D0),
				.a1(P05E0),
				.a2(P05F0),
				.a3(P06D0),
				.a4(P06E0),
				.a5(P06F0),
				.a6(P07D0),
				.a7(P07E0),
				.a8(P07F0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c005D2)
);

ninexnine_unit ninexnine_unit_1426(
				.clk(clk),
				.rstn(rstn),
				.a0(P05D1),
				.a1(P05E1),
				.a2(P05F1),
				.a3(P06D1),
				.a4(P06E1),
				.a5(P06F1),
				.a6(P07D1),
				.a7(P07E1),
				.a8(P07F1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c015D2)
);

ninexnine_unit ninexnine_unit_1427(
				.clk(clk),
				.rstn(rstn),
				.a0(P05D2),
				.a1(P05E2),
				.a2(P05F2),
				.a3(P06D2),
				.a4(P06E2),
				.a5(P06F2),
				.a6(P07D2),
				.a7(P07E2),
				.a8(P07F2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c025D2)
);

assign C05D2=c005D2+c015D2+c025D2;
assign A05D2=(C05D2>=0)?1:0;

ninexnine_unit ninexnine_unit_1428(
				.clk(clk),
				.rstn(rstn),
				.a0(P0600),
				.a1(P0610),
				.a2(P0620),
				.a3(P0700),
				.a4(P0710),
				.a5(P0720),
				.a6(P0800),
				.a7(P0810),
				.a8(P0820),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00602)
);

ninexnine_unit ninexnine_unit_1429(
				.clk(clk),
				.rstn(rstn),
				.a0(P0601),
				.a1(P0611),
				.a2(P0621),
				.a3(P0701),
				.a4(P0711),
				.a5(P0721),
				.a6(P0801),
				.a7(P0811),
				.a8(P0821),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01602)
);

ninexnine_unit ninexnine_unit_1430(
				.clk(clk),
				.rstn(rstn),
				.a0(P0602),
				.a1(P0612),
				.a2(P0622),
				.a3(P0702),
				.a4(P0712),
				.a5(P0722),
				.a6(P0802),
				.a7(P0812),
				.a8(P0822),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02602)
);

assign C0602=c00602+c01602+c02602;
assign A0602=(C0602>=0)?1:0;

ninexnine_unit ninexnine_unit_1431(
				.clk(clk),
				.rstn(rstn),
				.a0(P0610),
				.a1(P0620),
				.a2(P0630),
				.a3(P0710),
				.a4(P0720),
				.a5(P0730),
				.a6(P0810),
				.a7(P0820),
				.a8(P0830),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00612)
);

ninexnine_unit ninexnine_unit_1432(
				.clk(clk),
				.rstn(rstn),
				.a0(P0611),
				.a1(P0621),
				.a2(P0631),
				.a3(P0711),
				.a4(P0721),
				.a5(P0731),
				.a6(P0811),
				.a7(P0821),
				.a8(P0831),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01612)
);

ninexnine_unit ninexnine_unit_1433(
				.clk(clk),
				.rstn(rstn),
				.a0(P0612),
				.a1(P0622),
				.a2(P0632),
				.a3(P0712),
				.a4(P0722),
				.a5(P0732),
				.a6(P0812),
				.a7(P0822),
				.a8(P0832),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02612)
);

assign C0612=c00612+c01612+c02612;
assign A0612=(C0612>=0)?1:0;

ninexnine_unit ninexnine_unit_1434(
				.clk(clk),
				.rstn(rstn),
				.a0(P0620),
				.a1(P0630),
				.a2(P0640),
				.a3(P0720),
				.a4(P0730),
				.a5(P0740),
				.a6(P0820),
				.a7(P0830),
				.a8(P0840),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00622)
);

ninexnine_unit ninexnine_unit_1435(
				.clk(clk),
				.rstn(rstn),
				.a0(P0621),
				.a1(P0631),
				.a2(P0641),
				.a3(P0721),
				.a4(P0731),
				.a5(P0741),
				.a6(P0821),
				.a7(P0831),
				.a8(P0841),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01622)
);

ninexnine_unit ninexnine_unit_1436(
				.clk(clk),
				.rstn(rstn),
				.a0(P0622),
				.a1(P0632),
				.a2(P0642),
				.a3(P0722),
				.a4(P0732),
				.a5(P0742),
				.a6(P0822),
				.a7(P0832),
				.a8(P0842),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02622)
);

assign C0622=c00622+c01622+c02622;
assign A0622=(C0622>=0)?1:0;

ninexnine_unit ninexnine_unit_1437(
				.clk(clk),
				.rstn(rstn),
				.a0(P0630),
				.a1(P0640),
				.a2(P0650),
				.a3(P0730),
				.a4(P0740),
				.a5(P0750),
				.a6(P0830),
				.a7(P0840),
				.a8(P0850),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00632)
);

ninexnine_unit ninexnine_unit_1438(
				.clk(clk),
				.rstn(rstn),
				.a0(P0631),
				.a1(P0641),
				.a2(P0651),
				.a3(P0731),
				.a4(P0741),
				.a5(P0751),
				.a6(P0831),
				.a7(P0841),
				.a8(P0851),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01632)
);

ninexnine_unit ninexnine_unit_1439(
				.clk(clk),
				.rstn(rstn),
				.a0(P0632),
				.a1(P0642),
				.a2(P0652),
				.a3(P0732),
				.a4(P0742),
				.a5(P0752),
				.a6(P0832),
				.a7(P0842),
				.a8(P0852),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02632)
);

assign C0632=c00632+c01632+c02632;
assign A0632=(C0632>=0)?1:0;

ninexnine_unit ninexnine_unit_1440(
				.clk(clk),
				.rstn(rstn),
				.a0(P0640),
				.a1(P0650),
				.a2(P0660),
				.a3(P0740),
				.a4(P0750),
				.a5(P0760),
				.a6(P0840),
				.a7(P0850),
				.a8(P0860),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00642)
);

ninexnine_unit ninexnine_unit_1441(
				.clk(clk),
				.rstn(rstn),
				.a0(P0641),
				.a1(P0651),
				.a2(P0661),
				.a3(P0741),
				.a4(P0751),
				.a5(P0761),
				.a6(P0841),
				.a7(P0851),
				.a8(P0861),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01642)
);

ninexnine_unit ninexnine_unit_1442(
				.clk(clk),
				.rstn(rstn),
				.a0(P0642),
				.a1(P0652),
				.a2(P0662),
				.a3(P0742),
				.a4(P0752),
				.a5(P0762),
				.a6(P0842),
				.a7(P0852),
				.a8(P0862),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02642)
);

assign C0642=c00642+c01642+c02642;
assign A0642=(C0642>=0)?1:0;

ninexnine_unit ninexnine_unit_1443(
				.clk(clk),
				.rstn(rstn),
				.a0(P0650),
				.a1(P0660),
				.a2(P0670),
				.a3(P0750),
				.a4(P0760),
				.a5(P0770),
				.a6(P0850),
				.a7(P0860),
				.a8(P0870),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00652)
);

ninexnine_unit ninexnine_unit_1444(
				.clk(clk),
				.rstn(rstn),
				.a0(P0651),
				.a1(P0661),
				.a2(P0671),
				.a3(P0751),
				.a4(P0761),
				.a5(P0771),
				.a6(P0851),
				.a7(P0861),
				.a8(P0871),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01652)
);

ninexnine_unit ninexnine_unit_1445(
				.clk(clk),
				.rstn(rstn),
				.a0(P0652),
				.a1(P0662),
				.a2(P0672),
				.a3(P0752),
				.a4(P0762),
				.a5(P0772),
				.a6(P0852),
				.a7(P0862),
				.a8(P0872),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02652)
);

assign C0652=c00652+c01652+c02652;
assign A0652=(C0652>=0)?1:0;

ninexnine_unit ninexnine_unit_1446(
				.clk(clk),
				.rstn(rstn),
				.a0(P0660),
				.a1(P0670),
				.a2(P0680),
				.a3(P0760),
				.a4(P0770),
				.a5(P0780),
				.a6(P0860),
				.a7(P0870),
				.a8(P0880),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00662)
);

ninexnine_unit ninexnine_unit_1447(
				.clk(clk),
				.rstn(rstn),
				.a0(P0661),
				.a1(P0671),
				.a2(P0681),
				.a3(P0761),
				.a4(P0771),
				.a5(P0781),
				.a6(P0861),
				.a7(P0871),
				.a8(P0881),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01662)
);

ninexnine_unit ninexnine_unit_1448(
				.clk(clk),
				.rstn(rstn),
				.a0(P0662),
				.a1(P0672),
				.a2(P0682),
				.a3(P0762),
				.a4(P0772),
				.a5(P0782),
				.a6(P0862),
				.a7(P0872),
				.a8(P0882),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02662)
);

assign C0662=c00662+c01662+c02662;
assign A0662=(C0662>=0)?1:0;

ninexnine_unit ninexnine_unit_1449(
				.clk(clk),
				.rstn(rstn),
				.a0(P0670),
				.a1(P0680),
				.a2(P0690),
				.a3(P0770),
				.a4(P0780),
				.a5(P0790),
				.a6(P0870),
				.a7(P0880),
				.a8(P0890),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00672)
);

ninexnine_unit ninexnine_unit_1450(
				.clk(clk),
				.rstn(rstn),
				.a0(P0671),
				.a1(P0681),
				.a2(P0691),
				.a3(P0771),
				.a4(P0781),
				.a5(P0791),
				.a6(P0871),
				.a7(P0881),
				.a8(P0891),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01672)
);

ninexnine_unit ninexnine_unit_1451(
				.clk(clk),
				.rstn(rstn),
				.a0(P0672),
				.a1(P0682),
				.a2(P0692),
				.a3(P0772),
				.a4(P0782),
				.a5(P0792),
				.a6(P0872),
				.a7(P0882),
				.a8(P0892),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02672)
);

assign C0672=c00672+c01672+c02672;
assign A0672=(C0672>=0)?1:0;

ninexnine_unit ninexnine_unit_1452(
				.clk(clk),
				.rstn(rstn),
				.a0(P0680),
				.a1(P0690),
				.a2(P06A0),
				.a3(P0780),
				.a4(P0790),
				.a5(P07A0),
				.a6(P0880),
				.a7(P0890),
				.a8(P08A0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00682)
);

ninexnine_unit ninexnine_unit_1453(
				.clk(clk),
				.rstn(rstn),
				.a0(P0681),
				.a1(P0691),
				.a2(P06A1),
				.a3(P0781),
				.a4(P0791),
				.a5(P07A1),
				.a6(P0881),
				.a7(P0891),
				.a8(P08A1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01682)
);

ninexnine_unit ninexnine_unit_1454(
				.clk(clk),
				.rstn(rstn),
				.a0(P0682),
				.a1(P0692),
				.a2(P06A2),
				.a3(P0782),
				.a4(P0792),
				.a5(P07A2),
				.a6(P0882),
				.a7(P0892),
				.a8(P08A2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02682)
);

assign C0682=c00682+c01682+c02682;
assign A0682=(C0682>=0)?1:0;

ninexnine_unit ninexnine_unit_1455(
				.clk(clk),
				.rstn(rstn),
				.a0(P0690),
				.a1(P06A0),
				.a2(P06B0),
				.a3(P0790),
				.a4(P07A0),
				.a5(P07B0),
				.a6(P0890),
				.a7(P08A0),
				.a8(P08B0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00692)
);

ninexnine_unit ninexnine_unit_1456(
				.clk(clk),
				.rstn(rstn),
				.a0(P0691),
				.a1(P06A1),
				.a2(P06B1),
				.a3(P0791),
				.a4(P07A1),
				.a5(P07B1),
				.a6(P0891),
				.a7(P08A1),
				.a8(P08B1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01692)
);

ninexnine_unit ninexnine_unit_1457(
				.clk(clk),
				.rstn(rstn),
				.a0(P0692),
				.a1(P06A2),
				.a2(P06B2),
				.a3(P0792),
				.a4(P07A2),
				.a5(P07B2),
				.a6(P0892),
				.a7(P08A2),
				.a8(P08B2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02692)
);

assign C0692=c00692+c01692+c02692;
assign A0692=(C0692>=0)?1:0;

ninexnine_unit ninexnine_unit_1458(
				.clk(clk),
				.rstn(rstn),
				.a0(P06A0),
				.a1(P06B0),
				.a2(P06C0),
				.a3(P07A0),
				.a4(P07B0),
				.a5(P07C0),
				.a6(P08A0),
				.a7(P08B0),
				.a8(P08C0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c006A2)
);

ninexnine_unit ninexnine_unit_1459(
				.clk(clk),
				.rstn(rstn),
				.a0(P06A1),
				.a1(P06B1),
				.a2(P06C1),
				.a3(P07A1),
				.a4(P07B1),
				.a5(P07C1),
				.a6(P08A1),
				.a7(P08B1),
				.a8(P08C1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c016A2)
);

ninexnine_unit ninexnine_unit_1460(
				.clk(clk),
				.rstn(rstn),
				.a0(P06A2),
				.a1(P06B2),
				.a2(P06C2),
				.a3(P07A2),
				.a4(P07B2),
				.a5(P07C2),
				.a6(P08A2),
				.a7(P08B2),
				.a8(P08C2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c026A2)
);

assign C06A2=c006A2+c016A2+c026A2;
assign A06A2=(C06A2>=0)?1:0;

ninexnine_unit ninexnine_unit_1461(
				.clk(clk),
				.rstn(rstn),
				.a0(P06B0),
				.a1(P06C0),
				.a2(P06D0),
				.a3(P07B0),
				.a4(P07C0),
				.a5(P07D0),
				.a6(P08B0),
				.a7(P08C0),
				.a8(P08D0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c006B2)
);

ninexnine_unit ninexnine_unit_1462(
				.clk(clk),
				.rstn(rstn),
				.a0(P06B1),
				.a1(P06C1),
				.a2(P06D1),
				.a3(P07B1),
				.a4(P07C1),
				.a5(P07D1),
				.a6(P08B1),
				.a7(P08C1),
				.a8(P08D1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c016B2)
);

ninexnine_unit ninexnine_unit_1463(
				.clk(clk),
				.rstn(rstn),
				.a0(P06B2),
				.a1(P06C2),
				.a2(P06D2),
				.a3(P07B2),
				.a4(P07C2),
				.a5(P07D2),
				.a6(P08B2),
				.a7(P08C2),
				.a8(P08D2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c026B2)
);

assign C06B2=c006B2+c016B2+c026B2;
assign A06B2=(C06B2>=0)?1:0;

ninexnine_unit ninexnine_unit_1464(
				.clk(clk),
				.rstn(rstn),
				.a0(P06C0),
				.a1(P06D0),
				.a2(P06E0),
				.a3(P07C0),
				.a4(P07D0),
				.a5(P07E0),
				.a6(P08C0),
				.a7(P08D0),
				.a8(P08E0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c006C2)
);

ninexnine_unit ninexnine_unit_1465(
				.clk(clk),
				.rstn(rstn),
				.a0(P06C1),
				.a1(P06D1),
				.a2(P06E1),
				.a3(P07C1),
				.a4(P07D1),
				.a5(P07E1),
				.a6(P08C1),
				.a7(P08D1),
				.a8(P08E1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c016C2)
);

ninexnine_unit ninexnine_unit_1466(
				.clk(clk),
				.rstn(rstn),
				.a0(P06C2),
				.a1(P06D2),
				.a2(P06E2),
				.a3(P07C2),
				.a4(P07D2),
				.a5(P07E2),
				.a6(P08C2),
				.a7(P08D2),
				.a8(P08E2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c026C2)
);

assign C06C2=c006C2+c016C2+c026C2;
assign A06C2=(C06C2>=0)?1:0;

ninexnine_unit ninexnine_unit_1467(
				.clk(clk),
				.rstn(rstn),
				.a0(P06D0),
				.a1(P06E0),
				.a2(P06F0),
				.a3(P07D0),
				.a4(P07E0),
				.a5(P07F0),
				.a6(P08D0),
				.a7(P08E0),
				.a8(P08F0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c006D2)
);

ninexnine_unit ninexnine_unit_1468(
				.clk(clk),
				.rstn(rstn),
				.a0(P06D1),
				.a1(P06E1),
				.a2(P06F1),
				.a3(P07D1),
				.a4(P07E1),
				.a5(P07F1),
				.a6(P08D1),
				.a7(P08E1),
				.a8(P08F1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c016D2)
);

ninexnine_unit ninexnine_unit_1469(
				.clk(clk),
				.rstn(rstn),
				.a0(P06D2),
				.a1(P06E2),
				.a2(P06F2),
				.a3(P07D2),
				.a4(P07E2),
				.a5(P07F2),
				.a6(P08D2),
				.a7(P08E2),
				.a8(P08F2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c026D2)
);

assign C06D2=c006D2+c016D2+c026D2;
assign A06D2=(C06D2>=0)?1:0;

ninexnine_unit ninexnine_unit_1470(
				.clk(clk),
				.rstn(rstn),
				.a0(P0700),
				.a1(P0710),
				.a2(P0720),
				.a3(P0800),
				.a4(P0810),
				.a5(P0820),
				.a6(P0900),
				.a7(P0910),
				.a8(P0920),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00702)
);

ninexnine_unit ninexnine_unit_1471(
				.clk(clk),
				.rstn(rstn),
				.a0(P0701),
				.a1(P0711),
				.a2(P0721),
				.a3(P0801),
				.a4(P0811),
				.a5(P0821),
				.a6(P0901),
				.a7(P0911),
				.a8(P0921),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01702)
);

ninexnine_unit ninexnine_unit_1472(
				.clk(clk),
				.rstn(rstn),
				.a0(P0702),
				.a1(P0712),
				.a2(P0722),
				.a3(P0802),
				.a4(P0812),
				.a5(P0822),
				.a6(P0902),
				.a7(P0912),
				.a8(P0922),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02702)
);

assign C0702=c00702+c01702+c02702;
assign A0702=(C0702>=0)?1:0;

ninexnine_unit ninexnine_unit_1473(
				.clk(clk),
				.rstn(rstn),
				.a0(P0710),
				.a1(P0720),
				.a2(P0730),
				.a3(P0810),
				.a4(P0820),
				.a5(P0830),
				.a6(P0910),
				.a7(P0920),
				.a8(P0930),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00712)
);

ninexnine_unit ninexnine_unit_1474(
				.clk(clk),
				.rstn(rstn),
				.a0(P0711),
				.a1(P0721),
				.a2(P0731),
				.a3(P0811),
				.a4(P0821),
				.a5(P0831),
				.a6(P0911),
				.a7(P0921),
				.a8(P0931),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01712)
);

ninexnine_unit ninexnine_unit_1475(
				.clk(clk),
				.rstn(rstn),
				.a0(P0712),
				.a1(P0722),
				.a2(P0732),
				.a3(P0812),
				.a4(P0822),
				.a5(P0832),
				.a6(P0912),
				.a7(P0922),
				.a8(P0932),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02712)
);

assign C0712=c00712+c01712+c02712;
assign A0712=(C0712>=0)?1:0;

ninexnine_unit ninexnine_unit_1476(
				.clk(clk),
				.rstn(rstn),
				.a0(P0720),
				.a1(P0730),
				.a2(P0740),
				.a3(P0820),
				.a4(P0830),
				.a5(P0840),
				.a6(P0920),
				.a7(P0930),
				.a8(P0940),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00722)
);

ninexnine_unit ninexnine_unit_1477(
				.clk(clk),
				.rstn(rstn),
				.a0(P0721),
				.a1(P0731),
				.a2(P0741),
				.a3(P0821),
				.a4(P0831),
				.a5(P0841),
				.a6(P0921),
				.a7(P0931),
				.a8(P0941),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01722)
);

ninexnine_unit ninexnine_unit_1478(
				.clk(clk),
				.rstn(rstn),
				.a0(P0722),
				.a1(P0732),
				.a2(P0742),
				.a3(P0822),
				.a4(P0832),
				.a5(P0842),
				.a6(P0922),
				.a7(P0932),
				.a8(P0942),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02722)
);

assign C0722=c00722+c01722+c02722;
assign A0722=(C0722>=0)?1:0;

ninexnine_unit ninexnine_unit_1479(
				.clk(clk),
				.rstn(rstn),
				.a0(P0730),
				.a1(P0740),
				.a2(P0750),
				.a3(P0830),
				.a4(P0840),
				.a5(P0850),
				.a6(P0930),
				.a7(P0940),
				.a8(P0950),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00732)
);

ninexnine_unit ninexnine_unit_1480(
				.clk(clk),
				.rstn(rstn),
				.a0(P0731),
				.a1(P0741),
				.a2(P0751),
				.a3(P0831),
				.a4(P0841),
				.a5(P0851),
				.a6(P0931),
				.a7(P0941),
				.a8(P0951),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01732)
);

ninexnine_unit ninexnine_unit_1481(
				.clk(clk),
				.rstn(rstn),
				.a0(P0732),
				.a1(P0742),
				.a2(P0752),
				.a3(P0832),
				.a4(P0842),
				.a5(P0852),
				.a6(P0932),
				.a7(P0942),
				.a8(P0952),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02732)
);

assign C0732=c00732+c01732+c02732;
assign A0732=(C0732>=0)?1:0;

ninexnine_unit ninexnine_unit_1482(
				.clk(clk),
				.rstn(rstn),
				.a0(P0740),
				.a1(P0750),
				.a2(P0760),
				.a3(P0840),
				.a4(P0850),
				.a5(P0860),
				.a6(P0940),
				.a7(P0950),
				.a8(P0960),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00742)
);

ninexnine_unit ninexnine_unit_1483(
				.clk(clk),
				.rstn(rstn),
				.a0(P0741),
				.a1(P0751),
				.a2(P0761),
				.a3(P0841),
				.a4(P0851),
				.a5(P0861),
				.a6(P0941),
				.a7(P0951),
				.a8(P0961),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01742)
);

ninexnine_unit ninexnine_unit_1484(
				.clk(clk),
				.rstn(rstn),
				.a0(P0742),
				.a1(P0752),
				.a2(P0762),
				.a3(P0842),
				.a4(P0852),
				.a5(P0862),
				.a6(P0942),
				.a7(P0952),
				.a8(P0962),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02742)
);

assign C0742=c00742+c01742+c02742;
assign A0742=(C0742>=0)?1:0;

ninexnine_unit ninexnine_unit_1485(
				.clk(clk),
				.rstn(rstn),
				.a0(P0750),
				.a1(P0760),
				.a2(P0770),
				.a3(P0850),
				.a4(P0860),
				.a5(P0870),
				.a6(P0950),
				.a7(P0960),
				.a8(P0970),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00752)
);

ninexnine_unit ninexnine_unit_1486(
				.clk(clk),
				.rstn(rstn),
				.a0(P0751),
				.a1(P0761),
				.a2(P0771),
				.a3(P0851),
				.a4(P0861),
				.a5(P0871),
				.a6(P0951),
				.a7(P0961),
				.a8(P0971),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01752)
);

ninexnine_unit ninexnine_unit_1487(
				.clk(clk),
				.rstn(rstn),
				.a0(P0752),
				.a1(P0762),
				.a2(P0772),
				.a3(P0852),
				.a4(P0862),
				.a5(P0872),
				.a6(P0952),
				.a7(P0962),
				.a8(P0972),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02752)
);

assign C0752=c00752+c01752+c02752;
assign A0752=(C0752>=0)?1:0;

ninexnine_unit ninexnine_unit_1488(
				.clk(clk),
				.rstn(rstn),
				.a0(P0760),
				.a1(P0770),
				.a2(P0780),
				.a3(P0860),
				.a4(P0870),
				.a5(P0880),
				.a6(P0960),
				.a7(P0970),
				.a8(P0980),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00762)
);

ninexnine_unit ninexnine_unit_1489(
				.clk(clk),
				.rstn(rstn),
				.a0(P0761),
				.a1(P0771),
				.a2(P0781),
				.a3(P0861),
				.a4(P0871),
				.a5(P0881),
				.a6(P0961),
				.a7(P0971),
				.a8(P0981),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01762)
);

ninexnine_unit ninexnine_unit_1490(
				.clk(clk),
				.rstn(rstn),
				.a0(P0762),
				.a1(P0772),
				.a2(P0782),
				.a3(P0862),
				.a4(P0872),
				.a5(P0882),
				.a6(P0962),
				.a7(P0972),
				.a8(P0982),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02762)
);

assign C0762=c00762+c01762+c02762;
assign A0762=(C0762>=0)?1:0;

ninexnine_unit ninexnine_unit_1491(
				.clk(clk),
				.rstn(rstn),
				.a0(P0770),
				.a1(P0780),
				.a2(P0790),
				.a3(P0870),
				.a4(P0880),
				.a5(P0890),
				.a6(P0970),
				.a7(P0980),
				.a8(P0990),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00772)
);

ninexnine_unit ninexnine_unit_1492(
				.clk(clk),
				.rstn(rstn),
				.a0(P0771),
				.a1(P0781),
				.a2(P0791),
				.a3(P0871),
				.a4(P0881),
				.a5(P0891),
				.a6(P0971),
				.a7(P0981),
				.a8(P0991),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01772)
);

ninexnine_unit ninexnine_unit_1493(
				.clk(clk),
				.rstn(rstn),
				.a0(P0772),
				.a1(P0782),
				.a2(P0792),
				.a3(P0872),
				.a4(P0882),
				.a5(P0892),
				.a6(P0972),
				.a7(P0982),
				.a8(P0992),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02772)
);

assign C0772=c00772+c01772+c02772;
assign A0772=(C0772>=0)?1:0;

ninexnine_unit ninexnine_unit_1494(
				.clk(clk),
				.rstn(rstn),
				.a0(P0780),
				.a1(P0790),
				.a2(P07A0),
				.a3(P0880),
				.a4(P0890),
				.a5(P08A0),
				.a6(P0980),
				.a7(P0990),
				.a8(P09A0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00782)
);

ninexnine_unit ninexnine_unit_1495(
				.clk(clk),
				.rstn(rstn),
				.a0(P0781),
				.a1(P0791),
				.a2(P07A1),
				.a3(P0881),
				.a4(P0891),
				.a5(P08A1),
				.a6(P0981),
				.a7(P0991),
				.a8(P09A1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01782)
);

ninexnine_unit ninexnine_unit_1496(
				.clk(clk),
				.rstn(rstn),
				.a0(P0782),
				.a1(P0792),
				.a2(P07A2),
				.a3(P0882),
				.a4(P0892),
				.a5(P08A2),
				.a6(P0982),
				.a7(P0992),
				.a8(P09A2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02782)
);

assign C0782=c00782+c01782+c02782;
assign A0782=(C0782>=0)?1:0;

ninexnine_unit ninexnine_unit_1497(
				.clk(clk),
				.rstn(rstn),
				.a0(P0790),
				.a1(P07A0),
				.a2(P07B0),
				.a3(P0890),
				.a4(P08A0),
				.a5(P08B0),
				.a6(P0990),
				.a7(P09A0),
				.a8(P09B0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00792)
);

ninexnine_unit ninexnine_unit_1498(
				.clk(clk),
				.rstn(rstn),
				.a0(P0791),
				.a1(P07A1),
				.a2(P07B1),
				.a3(P0891),
				.a4(P08A1),
				.a5(P08B1),
				.a6(P0991),
				.a7(P09A1),
				.a8(P09B1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01792)
);

ninexnine_unit ninexnine_unit_1499(
				.clk(clk),
				.rstn(rstn),
				.a0(P0792),
				.a1(P07A2),
				.a2(P07B2),
				.a3(P0892),
				.a4(P08A2),
				.a5(P08B2),
				.a6(P0992),
				.a7(P09A2),
				.a8(P09B2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02792)
);

assign C0792=c00792+c01792+c02792;
assign A0792=(C0792>=0)?1:0;

ninexnine_unit ninexnine_unit_1500(
				.clk(clk),
				.rstn(rstn),
				.a0(P07A0),
				.a1(P07B0),
				.a2(P07C0),
				.a3(P08A0),
				.a4(P08B0),
				.a5(P08C0),
				.a6(P09A0),
				.a7(P09B0),
				.a8(P09C0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c007A2)
);

ninexnine_unit ninexnine_unit_1501(
				.clk(clk),
				.rstn(rstn),
				.a0(P07A1),
				.a1(P07B1),
				.a2(P07C1),
				.a3(P08A1),
				.a4(P08B1),
				.a5(P08C1),
				.a6(P09A1),
				.a7(P09B1),
				.a8(P09C1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c017A2)
);

ninexnine_unit ninexnine_unit_1502(
				.clk(clk),
				.rstn(rstn),
				.a0(P07A2),
				.a1(P07B2),
				.a2(P07C2),
				.a3(P08A2),
				.a4(P08B2),
				.a5(P08C2),
				.a6(P09A2),
				.a7(P09B2),
				.a8(P09C2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c027A2)
);

assign C07A2=c007A2+c017A2+c027A2;
assign A07A2=(C07A2>=0)?1:0;

ninexnine_unit ninexnine_unit_1503(
				.clk(clk),
				.rstn(rstn),
				.a0(P07B0),
				.a1(P07C0),
				.a2(P07D0),
				.a3(P08B0),
				.a4(P08C0),
				.a5(P08D0),
				.a6(P09B0),
				.a7(P09C0),
				.a8(P09D0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c007B2)
);

ninexnine_unit ninexnine_unit_1504(
				.clk(clk),
				.rstn(rstn),
				.a0(P07B1),
				.a1(P07C1),
				.a2(P07D1),
				.a3(P08B1),
				.a4(P08C1),
				.a5(P08D1),
				.a6(P09B1),
				.a7(P09C1),
				.a8(P09D1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c017B2)
);

ninexnine_unit ninexnine_unit_1505(
				.clk(clk),
				.rstn(rstn),
				.a0(P07B2),
				.a1(P07C2),
				.a2(P07D2),
				.a3(P08B2),
				.a4(P08C2),
				.a5(P08D2),
				.a6(P09B2),
				.a7(P09C2),
				.a8(P09D2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c027B2)
);

assign C07B2=c007B2+c017B2+c027B2;
assign A07B2=(C07B2>=0)?1:0;

ninexnine_unit ninexnine_unit_1506(
				.clk(clk),
				.rstn(rstn),
				.a0(P07C0),
				.a1(P07D0),
				.a2(P07E0),
				.a3(P08C0),
				.a4(P08D0),
				.a5(P08E0),
				.a6(P09C0),
				.a7(P09D0),
				.a8(P09E0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c007C2)
);

ninexnine_unit ninexnine_unit_1507(
				.clk(clk),
				.rstn(rstn),
				.a0(P07C1),
				.a1(P07D1),
				.a2(P07E1),
				.a3(P08C1),
				.a4(P08D1),
				.a5(P08E1),
				.a6(P09C1),
				.a7(P09D1),
				.a8(P09E1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c017C2)
);

ninexnine_unit ninexnine_unit_1508(
				.clk(clk),
				.rstn(rstn),
				.a0(P07C2),
				.a1(P07D2),
				.a2(P07E2),
				.a3(P08C2),
				.a4(P08D2),
				.a5(P08E2),
				.a6(P09C2),
				.a7(P09D2),
				.a8(P09E2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c027C2)
);

assign C07C2=c007C2+c017C2+c027C2;
assign A07C2=(C07C2>=0)?1:0;

ninexnine_unit ninexnine_unit_1509(
				.clk(clk),
				.rstn(rstn),
				.a0(P07D0),
				.a1(P07E0),
				.a2(P07F0),
				.a3(P08D0),
				.a4(P08E0),
				.a5(P08F0),
				.a6(P09D0),
				.a7(P09E0),
				.a8(P09F0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c007D2)
);

ninexnine_unit ninexnine_unit_1510(
				.clk(clk),
				.rstn(rstn),
				.a0(P07D1),
				.a1(P07E1),
				.a2(P07F1),
				.a3(P08D1),
				.a4(P08E1),
				.a5(P08F1),
				.a6(P09D1),
				.a7(P09E1),
				.a8(P09F1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c017D2)
);

ninexnine_unit ninexnine_unit_1511(
				.clk(clk),
				.rstn(rstn),
				.a0(P07D2),
				.a1(P07E2),
				.a2(P07F2),
				.a3(P08D2),
				.a4(P08E2),
				.a5(P08F2),
				.a6(P09D2),
				.a7(P09E2),
				.a8(P09F2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c027D2)
);

assign C07D2=c007D2+c017D2+c027D2;
assign A07D2=(C07D2>=0)?1:0;

ninexnine_unit ninexnine_unit_1512(
				.clk(clk),
				.rstn(rstn),
				.a0(P0800),
				.a1(P0810),
				.a2(P0820),
				.a3(P0900),
				.a4(P0910),
				.a5(P0920),
				.a6(P0A00),
				.a7(P0A10),
				.a8(P0A20),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00802)
);

ninexnine_unit ninexnine_unit_1513(
				.clk(clk),
				.rstn(rstn),
				.a0(P0801),
				.a1(P0811),
				.a2(P0821),
				.a3(P0901),
				.a4(P0911),
				.a5(P0921),
				.a6(P0A01),
				.a7(P0A11),
				.a8(P0A21),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01802)
);

ninexnine_unit ninexnine_unit_1514(
				.clk(clk),
				.rstn(rstn),
				.a0(P0802),
				.a1(P0812),
				.a2(P0822),
				.a3(P0902),
				.a4(P0912),
				.a5(P0922),
				.a6(P0A02),
				.a7(P0A12),
				.a8(P0A22),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02802)
);

assign C0802=c00802+c01802+c02802;
assign A0802=(C0802>=0)?1:0;

ninexnine_unit ninexnine_unit_1515(
				.clk(clk),
				.rstn(rstn),
				.a0(P0810),
				.a1(P0820),
				.a2(P0830),
				.a3(P0910),
				.a4(P0920),
				.a5(P0930),
				.a6(P0A10),
				.a7(P0A20),
				.a8(P0A30),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00812)
);

ninexnine_unit ninexnine_unit_1516(
				.clk(clk),
				.rstn(rstn),
				.a0(P0811),
				.a1(P0821),
				.a2(P0831),
				.a3(P0911),
				.a4(P0921),
				.a5(P0931),
				.a6(P0A11),
				.a7(P0A21),
				.a8(P0A31),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01812)
);

ninexnine_unit ninexnine_unit_1517(
				.clk(clk),
				.rstn(rstn),
				.a0(P0812),
				.a1(P0822),
				.a2(P0832),
				.a3(P0912),
				.a4(P0922),
				.a5(P0932),
				.a6(P0A12),
				.a7(P0A22),
				.a8(P0A32),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02812)
);

assign C0812=c00812+c01812+c02812;
assign A0812=(C0812>=0)?1:0;

ninexnine_unit ninexnine_unit_1518(
				.clk(clk),
				.rstn(rstn),
				.a0(P0820),
				.a1(P0830),
				.a2(P0840),
				.a3(P0920),
				.a4(P0930),
				.a5(P0940),
				.a6(P0A20),
				.a7(P0A30),
				.a8(P0A40),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00822)
);

ninexnine_unit ninexnine_unit_1519(
				.clk(clk),
				.rstn(rstn),
				.a0(P0821),
				.a1(P0831),
				.a2(P0841),
				.a3(P0921),
				.a4(P0931),
				.a5(P0941),
				.a6(P0A21),
				.a7(P0A31),
				.a8(P0A41),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01822)
);

ninexnine_unit ninexnine_unit_1520(
				.clk(clk),
				.rstn(rstn),
				.a0(P0822),
				.a1(P0832),
				.a2(P0842),
				.a3(P0922),
				.a4(P0932),
				.a5(P0942),
				.a6(P0A22),
				.a7(P0A32),
				.a8(P0A42),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02822)
);

assign C0822=c00822+c01822+c02822;
assign A0822=(C0822>=0)?1:0;

ninexnine_unit ninexnine_unit_1521(
				.clk(clk),
				.rstn(rstn),
				.a0(P0830),
				.a1(P0840),
				.a2(P0850),
				.a3(P0930),
				.a4(P0940),
				.a5(P0950),
				.a6(P0A30),
				.a7(P0A40),
				.a8(P0A50),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00832)
);

ninexnine_unit ninexnine_unit_1522(
				.clk(clk),
				.rstn(rstn),
				.a0(P0831),
				.a1(P0841),
				.a2(P0851),
				.a3(P0931),
				.a4(P0941),
				.a5(P0951),
				.a6(P0A31),
				.a7(P0A41),
				.a8(P0A51),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01832)
);

ninexnine_unit ninexnine_unit_1523(
				.clk(clk),
				.rstn(rstn),
				.a0(P0832),
				.a1(P0842),
				.a2(P0852),
				.a3(P0932),
				.a4(P0942),
				.a5(P0952),
				.a6(P0A32),
				.a7(P0A42),
				.a8(P0A52),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02832)
);

assign C0832=c00832+c01832+c02832;
assign A0832=(C0832>=0)?1:0;

ninexnine_unit ninexnine_unit_1524(
				.clk(clk),
				.rstn(rstn),
				.a0(P0840),
				.a1(P0850),
				.a2(P0860),
				.a3(P0940),
				.a4(P0950),
				.a5(P0960),
				.a6(P0A40),
				.a7(P0A50),
				.a8(P0A60),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00842)
);

ninexnine_unit ninexnine_unit_1525(
				.clk(clk),
				.rstn(rstn),
				.a0(P0841),
				.a1(P0851),
				.a2(P0861),
				.a3(P0941),
				.a4(P0951),
				.a5(P0961),
				.a6(P0A41),
				.a7(P0A51),
				.a8(P0A61),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01842)
);

ninexnine_unit ninexnine_unit_1526(
				.clk(clk),
				.rstn(rstn),
				.a0(P0842),
				.a1(P0852),
				.a2(P0862),
				.a3(P0942),
				.a4(P0952),
				.a5(P0962),
				.a6(P0A42),
				.a7(P0A52),
				.a8(P0A62),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02842)
);

assign C0842=c00842+c01842+c02842;
assign A0842=(C0842>=0)?1:0;

ninexnine_unit ninexnine_unit_1527(
				.clk(clk),
				.rstn(rstn),
				.a0(P0850),
				.a1(P0860),
				.a2(P0870),
				.a3(P0950),
				.a4(P0960),
				.a5(P0970),
				.a6(P0A50),
				.a7(P0A60),
				.a8(P0A70),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00852)
);

ninexnine_unit ninexnine_unit_1528(
				.clk(clk),
				.rstn(rstn),
				.a0(P0851),
				.a1(P0861),
				.a2(P0871),
				.a3(P0951),
				.a4(P0961),
				.a5(P0971),
				.a6(P0A51),
				.a7(P0A61),
				.a8(P0A71),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01852)
);

ninexnine_unit ninexnine_unit_1529(
				.clk(clk),
				.rstn(rstn),
				.a0(P0852),
				.a1(P0862),
				.a2(P0872),
				.a3(P0952),
				.a4(P0962),
				.a5(P0972),
				.a6(P0A52),
				.a7(P0A62),
				.a8(P0A72),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02852)
);

assign C0852=c00852+c01852+c02852;
assign A0852=(C0852>=0)?1:0;

ninexnine_unit ninexnine_unit_1530(
				.clk(clk),
				.rstn(rstn),
				.a0(P0860),
				.a1(P0870),
				.a2(P0880),
				.a3(P0960),
				.a4(P0970),
				.a5(P0980),
				.a6(P0A60),
				.a7(P0A70),
				.a8(P0A80),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00862)
);

ninexnine_unit ninexnine_unit_1531(
				.clk(clk),
				.rstn(rstn),
				.a0(P0861),
				.a1(P0871),
				.a2(P0881),
				.a3(P0961),
				.a4(P0971),
				.a5(P0981),
				.a6(P0A61),
				.a7(P0A71),
				.a8(P0A81),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01862)
);

ninexnine_unit ninexnine_unit_1532(
				.clk(clk),
				.rstn(rstn),
				.a0(P0862),
				.a1(P0872),
				.a2(P0882),
				.a3(P0962),
				.a4(P0972),
				.a5(P0982),
				.a6(P0A62),
				.a7(P0A72),
				.a8(P0A82),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02862)
);

assign C0862=c00862+c01862+c02862;
assign A0862=(C0862>=0)?1:0;

ninexnine_unit ninexnine_unit_1533(
				.clk(clk),
				.rstn(rstn),
				.a0(P0870),
				.a1(P0880),
				.a2(P0890),
				.a3(P0970),
				.a4(P0980),
				.a5(P0990),
				.a6(P0A70),
				.a7(P0A80),
				.a8(P0A90),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00872)
);

ninexnine_unit ninexnine_unit_1534(
				.clk(clk),
				.rstn(rstn),
				.a0(P0871),
				.a1(P0881),
				.a2(P0891),
				.a3(P0971),
				.a4(P0981),
				.a5(P0991),
				.a6(P0A71),
				.a7(P0A81),
				.a8(P0A91),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01872)
);

ninexnine_unit ninexnine_unit_1535(
				.clk(clk),
				.rstn(rstn),
				.a0(P0872),
				.a1(P0882),
				.a2(P0892),
				.a3(P0972),
				.a4(P0982),
				.a5(P0992),
				.a6(P0A72),
				.a7(P0A82),
				.a8(P0A92),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02872)
);

assign C0872=c00872+c01872+c02872;
assign A0872=(C0872>=0)?1:0;

ninexnine_unit ninexnine_unit_1536(
				.clk(clk),
				.rstn(rstn),
				.a0(P0880),
				.a1(P0890),
				.a2(P08A0),
				.a3(P0980),
				.a4(P0990),
				.a5(P09A0),
				.a6(P0A80),
				.a7(P0A90),
				.a8(P0AA0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00882)
);

ninexnine_unit ninexnine_unit_1537(
				.clk(clk),
				.rstn(rstn),
				.a0(P0881),
				.a1(P0891),
				.a2(P08A1),
				.a3(P0981),
				.a4(P0991),
				.a5(P09A1),
				.a6(P0A81),
				.a7(P0A91),
				.a8(P0AA1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01882)
);

ninexnine_unit ninexnine_unit_1538(
				.clk(clk),
				.rstn(rstn),
				.a0(P0882),
				.a1(P0892),
				.a2(P08A2),
				.a3(P0982),
				.a4(P0992),
				.a5(P09A2),
				.a6(P0A82),
				.a7(P0A92),
				.a8(P0AA2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02882)
);

assign C0882=c00882+c01882+c02882;
assign A0882=(C0882>=0)?1:0;

ninexnine_unit ninexnine_unit_1539(
				.clk(clk),
				.rstn(rstn),
				.a0(P0890),
				.a1(P08A0),
				.a2(P08B0),
				.a3(P0990),
				.a4(P09A0),
				.a5(P09B0),
				.a6(P0A90),
				.a7(P0AA0),
				.a8(P0AB0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00892)
);

ninexnine_unit ninexnine_unit_1540(
				.clk(clk),
				.rstn(rstn),
				.a0(P0891),
				.a1(P08A1),
				.a2(P08B1),
				.a3(P0991),
				.a4(P09A1),
				.a5(P09B1),
				.a6(P0A91),
				.a7(P0AA1),
				.a8(P0AB1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01892)
);

ninexnine_unit ninexnine_unit_1541(
				.clk(clk),
				.rstn(rstn),
				.a0(P0892),
				.a1(P08A2),
				.a2(P08B2),
				.a3(P0992),
				.a4(P09A2),
				.a5(P09B2),
				.a6(P0A92),
				.a7(P0AA2),
				.a8(P0AB2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02892)
);

assign C0892=c00892+c01892+c02892;
assign A0892=(C0892>=0)?1:0;

ninexnine_unit ninexnine_unit_1542(
				.clk(clk),
				.rstn(rstn),
				.a0(P08A0),
				.a1(P08B0),
				.a2(P08C0),
				.a3(P09A0),
				.a4(P09B0),
				.a5(P09C0),
				.a6(P0AA0),
				.a7(P0AB0),
				.a8(P0AC0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c008A2)
);

ninexnine_unit ninexnine_unit_1543(
				.clk(clk),
				.rstn(rstn),
				.a0(P08A1),
				.a1(P08B1),
				.a2(P08C1),
				.a3(P09A1),
				.a4(P09B1),
				.a5(P09C1),
				.a6(P0AA1),
				.a7(P0AB1),
				.a8(P0AC1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c018A2)
);

ninexnine_unit ninexnine_unit_1544(
				.clk(clk),
				.rstn(rstn),
				.a0(P08A2),
				.a1(P08B2),
				.a2(P08C2),
				.a3(P09A2),
				.a4(P09B2),
				.a5(P09C2),
				.a6(P0AA2),
				.a7(P0AB2),
				.a8(P0AC2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c028A2)
);

assign C08A2=c008A2+c018A2+c028A2;
assign A08A2=(C08A2>=0)?1:0;

ninexnine_unit ninexnine_unit_1545(
				.clk(clk),
				.rstn(rstn),
				.a0(P08B0),
				.a1(P08C0),
				.a2(P08D0),
				.a3(P09B0),
				.a4(P09C0),
				.a5(P09D0),
				.a6(P0AB0),
				.a7(P0AC0),
				.a8(P0AD0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c008B2)
);

ninexnine_unit ninexnine_unit_1546(
				.clk(clk),
				.rstn(rstn),
				.a0(P08B1),
				.a1(P08C1),
				.a2(P08D1),
				.a3(P09B1),
				.a4(P09C1),
				.a5(P09D1),
				.a6(P0AB1),
				.a7(P0AC1),
				.a8(P0AD1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c018B2)
);

ninexnine_unit ninexnine_unit_1547(
				.clk(clk),
				.rstn(rstn),
				.a0(P08B2),
				.a1(P08C2),
				.a2(P08D2),
				.a3(P09B2),
				.a4(P09C2),
				.a5(P09D2),
				.a6(P0AB2),
				.a7(P0AC2),
				.a8(P0AD2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c028B2)
);

assign C08B2=c008B2+c018B2+c028B2;
assign A08B2=(C08B2>=0)?1:0;

ninexnine_unit ninexnine_unit_1548(
				.clk(clk),
				.rstn(rstn),
				.a0(P08C0),
				.a1(P08D0),
				.a2(P08E0),
				.a3(P09C0),
				.a4(P09D0),
				.a5(P09E0),
				.a6(P0AC0),
				.a7(P0AD0),
				.a8(P0AE0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c008C2)
);

ninexnine_unit ninexnine_unit_1549(
				.clk(clk),
				.rstn(rstn),
				.a0(P08C1),
				.a1(P08D1),
				.a2(P08E1),
				.a3(P09C1),
				.a4(P09D1),
				.a5(P09E1),
				.a6(P0AC1),
				.a7(P0AD1),
				.a8(P0AE1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c018C2)
);

ninexnine_unit ninexnine_unit_1550(
				.clk(clk),
				.rstn(rstn),
				.a0(P08C2),
				.a1(P08D2),
				.a2(P08E2),
				.a3(P09C2),
				.a4(P09D2),
				.a5(P09E2),
				.a6(P0AC2),
				.a7(P0AD2),
				.a8(P0AE2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c028C2)
);

assign C08C2=c008C2+c018C2+c028C2;
assign A08C2=(C08C2>=0)?1:0;

ninexnine_unit ninexnine_unit_1551(
				.clk(clk),
				.rstn(rstn),
				.a0(P08D0),
				.a1(P08E0),
				.a2(P08F0),
				.a3(P09D0),
				.a4(P09E0),
				.a5(P09F0),
				.a6(P0AD0),
				.a7(P0AE0),
				.a8(P0AF0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c008D2)
);

ninexnine_unit ninexnine_unit_1552(
				.clk(clk),
				.rstn(rstn),
				.a0(P08D1),
				.a1(P08E1),
				.a2(P08F1),
				.a3(P09D1),
				.a4(P09E1),
				.a5(P09F1),
				.a6(P0AD1),
				.a7(P0AE1),
				.a8(P0AF1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c018D2)
);

ninexnine_unit ninexnine_unit_1553(
				.clk(clk),
				.rstn(rstn),
				.a0(P08D2),
				.a1(P08E2),
				.a2(P08F2),
				.a3(P09D2),
				.a4(P09E2),
				.a5(P09F2),
				.a6(P0AD2),
				.a7(P0AE2),
				.a8(P0AF2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c028D2)
);

assign C08D2=c008D2+c018D2+c028D2;
assign A08D2=(C08D2>=0)?1:0;

ninexnine_unit ninexnine_unit_1554(
				.clk(clk),
				.rstn(rstn),
				.a0(P0900),
				.a1(P0910),
				.a2(P0920),
				.a3(P0A00),
				.a4(P0A10),
				.a5(P0A20),
				.a6(P0B00),
				.a7(P0B10),
				.a8(P0B20),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00902)
);

ninexnine_unit ninexnine_unit_1555(
				.clk(clk),
				.rstn(rstn),
				.a0(P0901),
				.a1(P0911),
				.a2(P0921),
				.a3(P0A01),
				.a4(P0A11),
				.a5(P0A21),
				.a6(P0B01),
				.a7(P0B11),
				.a8(P0B21),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01902)
);

ninexnine_unit ninexnine_unit_1556(
				.clk(clk),
				.rstn(rstn),
				.a0(P0902),
				.a1(P0912),
				.a2(P0922),
				.a3(P0A02),
				.a4(P0A12),
				.a5(P0A22),
				.a6(P0B02),
				.a7(P0B12),
				.a8(P0B22),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02902)
);

assign C0902=c00902+c01902+c02902;
assign A0902=(C0902>=0)?1:0;

ninexnine_unit ninexnine_unit_1557(
				.clk(clk),
				.rstn(rstn),
				.a0(P0910),
				.a1(P0920),
				.a2(P0930),
				.a3(P0A10),
				.a4(P0A20),
				.a5(P0A30),
				.a6(P0B10),
				.a7(P0B20),
				.a8(P0B30),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00912)
);

ninexnine_unit ninexnine_unit_1558(
				.clk(clk),
				.rstn(rstn),
				.a0(P0911),
				.a1(P0921),
				.a2(P0931),
				.a3(P0A11),
				.a4(P0A21),
				.a5(P0A31),
				.a6(P0B11),
				.a7(P0B21),
				.a8(P0B31),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01912)
);

ninexnine_unit ninexnine_unit_1559(
				.clk(clk),
				.rstn(rstn),
				.a0(P0912),
				.a1(P0922),
				.a2(P0932),
				.a3(P0A12),
				.a4(P0A22),
				.a5(P0A32),
				.a6(P0B12),
				.a7(P0B22),
				.a8(P0B32),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02912)
);

assign C0912=c00912+c01912+c02912;
assign A0912=(C0912>=0)?1:0;

ninexnine_unit ninexnine_unit_1560(
				.clk(clk),
				.rstn(rstn),
				.a0(P0920),
				.a1(P0930),
				.a2(P0940),
				.a3(P0A20),
				.a4(P0A30),
				.a5(P0A40),
				.a6(P0B20),
				.a7(P0B30),
				.a8(P0B40),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00922)
);

ninexnine_unit ninexnine_unit_1561(
				.clk(clk),
				.rstn(rstn),
				.a0(P0921),
				.a1(P0931),
				.a2(P0941),
				.a3(P0A21),
				.a4(P0A31),
				.a5(P0A41),
				.a6(P0B21),
				.a7(P0B31),
				.a8(P0B41),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01922)
);

ninexnine_unit ninexnine_unit_1562(
				.clk(clk),
				.rstn(rstn),
				.a0(P0922),
				.a1(P0932),
				.a2(P0942),
				.a3(P0A22),
				.a4(P0A32),
				.a5(P0A42),
				.a6(P0B22),
				.a7(P0B32),
				.a8(P0B42),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02922)
);

assign C0922=c00922+c01922+c02922;
assign A0922=(C0922>=0)?1:0;

ninexnine_unit ninexnine_unit_1563(
				.clk(clk),
				.rstn(rstn),
				.a0(P0930),
				.a1(P0940),
				.a2(P0950),
				.a3(P0A30),
				.a4(P0A40),
				.a5(P0A50),
				.a6(P0B30),
				.a7(P0B40),
				.a8(P0B50),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00932)
);

ninexnine_unit ninexnine_unit_1564(
				.clk(clk),
				.rstn(rstn),
				.a0(P0931),
				.a1(P0941),
				.a2(P0951),
				.a3(P0A31),
				.a4(P0A41),
				.a5(P0A51),
				.a6(P0B31),
				.a7(P0B41),
				.a8(P0B51),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01932)
);

ninexnine_unit ninexnine_unit_1565(
				.clk(clk),
				.rstn(rstn),
				.a0(P0932),
				.a1(P0942),
				.a2(P0952),
				.a3(P0A32),
				.a4(P0A42),
				.a5(P0A52),
				.a6(P0B32),
				.a7(P0B42),
				.a8(P0B52),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02932)
);

assign C0932=c00932+c01932+c02932;
assign A0932=(C0932>=0)?1:0;

ninexnine_unit ninexnine_unit_1566(
				.clk(clk),
				.rstn(rstn),
				.a0(P0940),
				.a1(P0950),
				.a2(P0960),
				.a3(P0A40),
				.a4(P0A50),
				.a5(P0A60),
				.a6(P0B40),
				.a7(P0B50),
				.a8(P0B60),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00942)
);

ninexnine_unit ninexnine_unit_1567(
				.clk(clk),
				.rstn(rstn),
				.a0(P0941),
				.a1(P0951),
				.a2(P0961),
				.a3(P0A41),
				.a4(P0A51),
				.a5(P0A61),
				.a6(P0B41),
				.a7(P0B51),
				.a8(P0B61),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01942)
);

ninexnine_unit ninexnine_unit_1568(
				.clk(clk),
				.rstn(rstn),
				.a0(P0942),
				.a1(P0952),
				.a2(P0962),
				.a3(P0A42),
				.a4(P0A52),
				.a5(P0A62),
				.a6(P0B42),
				.a7(P0B52),
				.a8(P0B62),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02942)
);

assign C0942=c00942+c01942+c02942;
assign A0942=(C0942>=0)?1:0;

ninexnine_unit ninexnine_unit_1569(
				.clk(clk),
				.rstn(rstn),
				.a0(P0950),
				.a1(P0960),
				.a2(P0970),
				.a3(P0A50),
				.a4(P0A60),
				.a5(P0A70),
				.a6(P0B50),
				.a7(P0B60),
				.a8(P0B70),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00952)
);

ninexnine_unit ninexnine_unit_1570(
				.clk(clk),
				.rstn(rstn),
				.a0(P0951),
				.a1(P0961),
				.a2(P0971),
				.a3(P0A51),
				.a4(P0A61),
				.a5(P0A71),
				.a6(P0B51),
				.a7(P0B61),
				.a8(P0B71),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01952)
);

ninexnine_unit ninexnine_unit_1571(
				.clk(clk),
				.rstn(rstn),
				.a0(P0952),
				.a1(P0962),
				.a2(P0972),
				.a3(P0A52),
				.a4(P0A62),
				.a5(P0A72),
				.a6(P0B52),
				.a7(P0B62),
				.a8(P0B72),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02952)
);

assign C0952=c00952+c01952+c02952;
assign A0952=(C0952>=0)?1:0;

ninexnine_unit ninexnine_unit_1572(
				.clk(clk),
				.rstn(rstn),
				.a0(P0960),
				.a1(P0970),
				.a2(P0980),
				.a3(P0A60),
				.a4(P0A70),
				.a5(P0A80),
				.a6(P0B60),
				.a7(P0B70),
				.a8(P0B80),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00962)
);

ninexnine_unit ninexnine_unit_1573(
				.clk(clk),
				.rstn(rstn),
				.a0(P0961),
				.a1(P0971),
				.a2(P0981),
				.a3(P0A61),
				.a4(P0A71),
				.a5(P0A81),
				.a6(P0B61),
				.a7(P0B71),
				.a8(P0B81),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01962)
);

ninexnine_unit ninexnine_unit_1574(
				.clk(clk),
				.rstn(rstn),
				.a0(P0962),
				.a1(P0972),
				.a2(P0982),
				.a3(P0A62),
				.a4(P0A72),
				.a5(P0A82),
				.a6(P0B62),
				.a7(P0B72),
				.a8(P0B82),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02962)
);

assign C0962=c00962+c01962+c02962;
assign A0962=(C0962>=0)?1:0;

ninexnine_unit ninexnine_unit_1575(
				.clk(clk),
				.rstn(rstn),
				.a0(P0970),
				.a1(P0980),
				.a2(P0990),
				.a3(P0A70),
				.a4(P0A80),
				.a5(P0A90),
				.a6(P0B70),
				.a7(P0B80),
				.a8(P0B90),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00972)
);

ninexnine_unit ninexnine_unit_1576(
				.clk(clk),
				.rstn(rstn),
				.a0(P0971),
				.a1(P0981),
				.a2(P0991),
				.a3(P0A71),
				.a4(P0A81),
				.a5(P0A91),
				.a6(P0B71),
				.a7(P0B81),
				.a8(P0B91),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01972)
);

ninexnine_unit ninexnine_unit_1577(
				.clk(clk),
				.rstn(rstn),
				.a0(P0972),
				.a1(P0982),
				.a2(P0992),
				.a3(P0A72),
				.a4(P0A82),
				.a5(P0A92),
				.a6(P0B72),
				.a7(P0B82),
				.a8(P0B92),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02972)
);

assign C0972=c00972+c01972+c02972;
assign A0972=(C0972>=0)?1:0;

ninexnine_unit ninexnine_unit_1578(
				.clk(clk),
				.rstn(rstn),
				.a0(P0980),
				.a1(P0990),
				.a2(P09A0),
				.a3(P0A80),
				.a4(P0A90),
				.a5(P0AA0),
				.a6(P0B80),
				.a7(P0B90),
				.a8(P0BA0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00982)
);

ninexnine_unit ninexnine_unit_1579(
				.clk(clk),
				.rstn(rstn),
				.a0(P0981),
				.a1(P0991),
				.a2(P09A1),
				.a3(P0A81),
				.a4(P0A91),
				.a5(P0AA1),
				.a6(P0B81),
				.a7(P0B91),
				.a8(P0BA1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01982)
);

ninexnine_unit ninexnine_unit_1580(
				.clk(clk),
				.rstn(rstn),
				.a0(P0982),
				.a1(P0992),
				.a2(P09A2),
				.a3(P0A82),
				.a4(P0A92),
				.a5(P0AA2),
				.a6(P0B82),
				.a7(P0B92),
				.a8(P0BA2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02982)
);

assign C0982=c00982+c01982+c02982;
assign A0982=(C0982>=0)?1:0;

ninexnine_unit ninexnine_unit_1581(
				.clk(clk),
				.rstn(rstn),
				.a0(P0990),
				.a1(P09A0),
				.a2(P09B0),
				.a3(P0A90),
				.a4(P0AA0),
				.a5(P0AB0),
				.a6(P0B90),
				.a7(P0BA0),
				.a8(P0BB0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00992)
);

ninexnine_unit ninexnine_unit_1582(
				.clk(clk),
				.rstn(rstn),
				.a0(P0991),
				.a1(P09A1),
				.a2(P09B1),
				.a3(P0A91),
				.a4(P0AA1),
				.a5(P0AB1),
				.a6(P0B91),
				.a7(P0BA1),
				.a8(P0BB1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01992)
);

ninexnine_unit ninexnine_unit_1583(
				.clk(clk),
				.rstn(rstn),
				.a0(P0992),
				.a1(P09A2),
				.a2(P09B2),
				.a3(P0A92),
				.a4(P0AA2),
				.a5(P0AB2),
				.a6(P0B92),
				.a7(P0BA2),
				.a8(P0BB2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02992)
);

assign C0992=c00992+c01992+c02992;
assign A0992=(C0992>=0)?1:0;

ninexnine_unit ninexnine_unit_1584(
				.clk(clk),
				.rstn(rstn),
				.a0(P09A0),
				.a1(P09B0),
				.a2(P09C0),
				.a3(P0AA0),
				.a4(P0AB0),
				.a5(P0AC0),
				.a6(P0BA0),
				.a7(P0BB0),
				.a8(P0BC0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c009A2)
);

ninexnine_unit ninexnine_unit_1585(
				.clk(clk),
				.rstn(rstn),
				.a0(P09A1),
				.a1(P09B1),
				.a2(P09C1),
				.a3(P0AA1),
				.a4(P0AB1),
				.a5(P0AC1),
				.a6(P0BA1),
				.a7(P0BB1),
				.a8(P0BC1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c019A2)
);

ninexnine_unit ninexnine_unit_1586(
				.clk(clk),
				.rstn(rstn),
				.a0(P09A2),
				.a1(P09B2),
				.a2(P09C2),
				.a3(P0AA2),
				.a4(P0AB2),
				.a5(P0AC2),
				.a6(P0BA2),
				.a7(P0BB2),
				.a8(P0BC2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c029A2)
);

assign C09A2=c009A2+c019A2+c029A2;
assign A09A2=(C09A2>=0)?1:0;

ninexnine_unit ninexnine_unit_1587(
				.clk(clk),
				.rstn(rstn),
				.a0(P09B0),
				.a1(P09C0),
				.a2(P09D0),
				.a3(P0AB0),
				.a4(P0AC0),
				.a5(P0AD0),
				.a6(P0BB0),
				.a7(P0BC0),
				.a8(P0BD0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c009B2)
);

ninexnine_unit ninexnine_unit_1588(
				.clk(clk),
				.rstn(rstn),
				.a0(P09B1),
				.a1(P09C1),
				.a2(P09D1),
				.a3(P0AB1),
				.a4(P0AC1),
				.a5(P0AD1),
				.a6(P0BB1),
				.a7(P0BC1),
				.a8(P0BD1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c019B2)
);

ninexnine_unit ninexnine_unit_1589(
				.clk(clk),
				.rstn(rstn),
				.a0(P09B2),
				.a1(P09C2),
				.a2(P09D2),
				.a3(P0AB2),
				.a4(P0AC2),
				.a5(P0AD2),
				.a6(P0BB2),
				.a7(P0BC2),
				.a8(P0BD2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c029B2)
);

assign C09B2=c009B2+c019B2+c029B2;
assign A09B2=(C09B2>=0)?1:0;

ninexnine_unit ninexnine_unit_1590(
				.clk(clk),
				.rstn(rstn),
				.a0(P09C0),
				.a1(P09D0),
				.a2(P09E0),
				.a3(P0AC0),
				.a4(P0AD0),
				.a5(P0AE0),
				.a6(P0BC0),
				.a7(P0BD0),
				.a8(P0BE0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c009C2)
);

ninexnine_unit ninexnine_unit_1591(
				.clk(clk),
				.rstn(rstn),
				.a0(P09C1),
				.a1(P09D1),
				.a2(P09E1),
				.a3(P0AC1),
				.a4(P0AD1),
				.a5(P0AE1),
				.a6(P0BC1),
				.a7(P0BD1),
				.a8(P0BE1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c019C2)
);

ninexnine_unit ninexnine_unit_1592(
				.clk(clk),
				.rstn(rstn),
				.a0(P09C2),
				.a1(P09D2),
				.a2(P09E2),
				.a3(P0AC2),
				.a4(P0AD2),
				.a5(P0AE2),
				.a6(P0BC2),
				.a7(P0BD2),
				.a8(P0BE2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c029C2)
);

assign C09C2=c009C2+c019C2+c029C2;
assign A09C2=(C09C2>=0)?1:0;

ninexnine_unit ninexnine_unit_1593(
				.clk(clk),
				.rstn(rstn),
				.a0(P09D0),
				.a1(P09E0),
				.a2(P09F0),
				.a3(P0AD0),
				.a4(P0AE0),
				.a5(P0AF0),
				.a6(P0BD0),
				.a7(P0BE0),
				.a8(P0BF0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c009D2)
);

ninexnine_unit ninexnine_unit_1594(
				.clk(clk),
				.rstn(rstn),
				.a0(P09D1),
				.a1(P09E1),
				.a2(P09F1),
				.a3(P0AD1),
				.a4(P0AE1),
				.a5(P0AF1),
				.a6(P0BD1),
				.a7(P0BE1),
				.a8(P0BF1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c019D2)
);

ninexnine_unit ninexnine_unit_1595(
				.clk(clk),
				.rstn(rstn),
				.a0(P09D2),
				.a1(P09E2),
				.a2(P09F2),
				.a3(P0AD2),
				.a4(P0AE2),
				.a5(P0AF2),
				.a6(P0BD2),
				.a7(P0BE2),
				.a8(P0BF2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c029D2)
);

assign C09D2=c009D2+c019D2+c029D2;
assign A09D2=(C09D2>=0)?1:0;

ninexnine_unit ninexnine_unit_1596(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A00),
				.a1(P0A10),
				.a2(P0A20),
				.a3(P0B00),
				.a4(P0B10),
				.a5(P0B20),
				.a6(P0C00),
				.a7(P0C10),
				.a8(P0C20),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00A02)
);

ninexnine_unit ninexnine_unit_1597(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A01),
				.a1(P0A11),
				.a2(P0A21),
				.a3(P0B01),
				.a4(P0B11),
				.a5(P0B21),
				.a6(P0C01),
				.a7(P0C11),
				.a8(P0C21),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01A02)
);

ninexnine_unit ninexnine_unit_1598(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A02),
				.a1(P0A12),
				.a2(P0A22),
				.a3(P0B02),
				.a4(P0B12),
				.a5(P0B22),
				.a6(P0C02),
				.a7(P0C12),
				.a8(P0C22),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02A02)
);

assign C0A02=c00A02+c01A02+c02A02;
assign A0A02=(C0A02>=0)?1:0;

ninexnine_unit ninexnine_unit_1599(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A10),
				.a1(P0A20),
				.a2(P0A30),
				.a3(P0B10),
				.a4(P0B20),
				.a5(P0B30),
				.a6(P0C10),
				.a7(P0C20),
				.a8(P0C30),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00A12)
);

ninexnine_unit ninexnine_unit_1600(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A11),
				.a1(P0A21),
				.a2(P0A31),
				.a3(P0B11),
				.a4(P0B21),
				.a5(P0B31),
				.a6(P0C11),
				.a7(P0C21),
				.a8(P0C31),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01A12)
);

ninexnine_unit ninexnine_unit_1601(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A12),
				.a1(P0A22),
				.a2(P0A32),
				.a3(P0B12),
				.a4(P0B22),
				.a5(P0B32),
				.a6(P0C12),
				.a7(P0C22),
				.a8(P0C32),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02A12)
);

assign C0A12=c00A12+c01A12+c02A12;
assign A0A12=(C0A12>=0)?1:0;

ninexnine_unit ninexnine_unit_1602(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A20),
				.a1(P0A30),
				.a2(P0A40),
				.a3(P0B20),
				.a4(P0B30),
				.a5(P0B40),
				.a6(P0C20),
				.a7(P0C30),
				.a8(P0C40),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00A22)
);

ninexnine_unit ninexnine_unit_1603(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A21),
				.a1(P0A31),
				.a2(P0A41),
				.a3(P0B21),
				.a4(P0B31),
				.a5(P0B41),
				.a6(P0C21),
				.a7(P0C31),
				.a8(P0C41),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01A22)
);

ninexnine_unit ninexnine_unit_1604(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A22),
				.a1(P0A32),
				.a2(P0A42),
				.a3(P0B22),
				.a4(P0B32),
				.a5(P0B42),
				.a6(P0C22),
				.a7(P0C32),
				.a8(P0C42),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02A22)
);

assign C0A22=c00A22+c01A22+c02A22;
assign A0A22=(C0A22>=0)?1:0;

ninexnine_unit ninexnine_unit_1605(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A30),
				.a1(P0A40),
				.a2(P0A50),
				.a3(P0B30),
				.a4(P0B40),
				.a5(P0B50),
				.a6(P0C30),
				.a7(P0C40),
				.a8(P0C50),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00A32)
);

ninexnine_unit ninexnine_unit_1606(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A31),
				.a1(P0A41),
				.a2(P0A51),
				.a3(P0B31),
				.a4(P0B41),
				.a5(P0B51),
				.a6(P0C31),
				.a7(P0C41),
				.a8(P0C51),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01A32)
);

ninexnine_unit ninexnine_unit_1607(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A32),
				.a1(P0A42),
				.a2(P0A52),
				.a3(P0B32),
				.a4(P0B42),
				.a5(P0B52),
				.a6(P0C32),
				.a7(P0C42),
				.a8(P0C52),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02A32)
);

assign C0A32=c00A32+c01A32+c02A32;
assign A0A32=(C0A32>=0)?1:0;

ninexnine_unit ninexnine_unit_1608(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A40),
				.a1(P0A50),
				.a2(P0A60),
				.a3(P0B40),
				.a4(P0B50),
				.a5(P0B60),
				.a6(P0C40),
				.a7(P0C50),
				.a8(P0C60),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00A42)
);

ninexnine_unit ninexnine_unit_1609(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A41),
				.a1(P0A51),
				.a2(P0A61),
				.a3(P0B41),
				.a4(P0B51),
				.a5(P0B61),
				.a6(P0C41),
				.a7(P0C51),
				.a8(P0C61),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01A42)
);

ninexnine_unit ninexnine_unit_1610(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A42),
				.a1(P0A52),
				.a2(P0A62),
				.a3(P0B42),
				.a4(P0B52),
				.a5(P0B62),
				.a6(P0C42),
				.a7(P0C52),
				.a8(P0C62),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02A42)
);

assign C0A42=c00A42+c01A42+c02A42;
assign A0A42=(C0A42>=0)?1:0;

ninexnine_unit ninexnine_unit_1611(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A50),
				.a1(P0A60),
				.a2(P0A70),
				.a3(P0B50),
				.a4(P0B60),
				.a5(P0B70),
				.a6(P0C50),
				.a7(P0C60),
				.a8(P0C70),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00A52)
);

ninexnine_unit ninexnine_unit_1612(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A51),
				.a1(P0A61),
				.a2(P0A71),
				.a3(P0B51),
				.a4(P0B61),
				.a5(P0B71),
				.a6(P0C51),
				.a7(P0C61),
				.a8(P0C71),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01A52)
);

ninexnine_unit ninexnine_unit_1613(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A52),
				.a1(P0A62),
				.a2(P0A72),
				.a3(P0B52),
				.a4(P0B62),
				.a5(P0B72),
				.a6(P0C52),
				.a7(P0C62),
				.a8(P0C72),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02A52)
);

assign C0A52=c00A52+c01A52+c02A52;
assign A0A52=(C0A52>=0)?1:0;

ninexnine_unit ninexnine_unit_1614(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A60),
				.a1(P0A70),
				.a2(P0A80),
				.a3(P0B60),
				.a4(P0B70),
				.a5(P0B80),
				.a6(P0C60),
				.a7(P0C70),
				.a8(P0C80),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00A62)
);

ninexnine_unit ninexnine_unit_1615(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A61),
				.a1(P0A71),
				.a2(P0A81),
				.a3(P0B61),
				.a4(P0B71),
				.a5(P0B81),
				.a6(P0C61),
				.a7(P0C71),
				.a8(P0C81),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01A62)
);

ninexnine_unit ninexnine_unit_1616(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A62),
				.a1(P0A72),
				.a2(P0A82),
				.a3(P0B62),
				.a4(P0B72),
				.a5(P0B82),
				.a6(P0C62),
				.a7(P0C72),
				.a8(P0C82),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02A62)
);

assign C0A62=c00A62+c01A62+c02A62;
assign A0A62=(C0A62>=0)?1:0;

ninexnine_unit ninexnine_unit_1617(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A70),
				.a1(P0A80),
				.a2(P0A90),
				.a3(P0B70),
				.a4(P0B80),
				.a5(P0B90),
				.a6(P0C70),
				.a7(P0C80),
				.a8(P0C90),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00A72)
);

ninexnine_unit ninexnine_unit_1618(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A71),
				.a1(P0A81),
				.a2(P0A91),
				.a3(P0B71),
				.a4(P0B81),
				.a5(P0B91),
				.a6(P0C71),
				.a7(P0C81),
				.a8(P0C91),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01A72)
);

ninexnine_unit ninexnine_unit_1619(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A72),
				.a1(P0A82),
				.a2(P0A92),
				.a3(P0B72),
				.a4(P0B82),
				.a5(P0B92),
				.a6(P0C72),
				.a7(P0C82),
				.a8(P0C92),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02A72)
);

assign C0A72=c00A72+c01A72+c02A72;
assign A0A72=(C0A72>=0)?1:0;

ninexnine_unit ninexnine_unit_1620(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A80),
				.a1(P0A90),
				.a2(P0AA0),
				.a3(P0B80),
				.a4(P0B90),
				.a5(P0BA0),
				.a6(P0C80),
				.a7(P0C90),
				.a8(P0CA0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00A82)
);

ninexnine_unit ninexnine_unit_1621(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A81),
				.a1(P0A91),
				.a2(P0AA1),
				.a3(P0B81),
				.a4(P0B91),
				.a5(P0BA1),
				.a6(P0C81),
				.a7(P0C91),
				.a8(P0CA1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01A82)
);

ninexnine_unit ninexnine_unit_1622(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A82),
				.a1(P0A92),
				.a2(P0AA2),
				.a3(P0B82),
				.a4(P0B92),
				.a5(P0BA2),
				.a6(P0C82),
				.a7(P0C92),
				.a8(P0CA2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02A82)
);

assign C0A82=c00A82+c01A82+c02A82;
assign A0A82=(C0A82>=0)?1:0;

ninexnine_unit ninexnine_unit_1623(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A90),
				.a1(P0AA0),
				.a2(P0AB0),
				.a3(P0B90),
				.a4(P0BA0),
				.a5(P0BB0),
				.a6(P0C90),
				.a7(P0CA0),
				.a8(P0CB0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00A92)
);

ninexnine_unit ninexnine_unit_1624(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A91),
				.a1(P0AA1),
				.a2(P0AB1),
				.a3(P0B91),
				.a4(P0BA1),
				.a5(P0BB1),
				.a6(P0C91),
				.a7(P0CA1),
				.a8(P0CB1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01A92)
);

ninexnine_unit ninexnine_unit_1625(
				.clk(clk),
				.rstn(rstn),
				.a0(P0A92),
				.a1(P0AA2),
				.a2(P0AB2),
				.a3(P0B92),
				.a4(P0BA2),
				.a5(P0BB2),
				.a6(P0C92),
				.a7(P0CA2),
				.a8(P0CB2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02A92)
);

assign C0A92=c00A92+c01A92+c02A92;
assign A0A92=(C0A92>=0)?1:0;

ninexnine_unit ninexnine_unit_1626(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AA0),
				.a1(P0AB0),
				.a2(P0AC0),
				.a3(P0BA0),
				.a4(P0BB0),
				.a5(P0BC0),
				.a6(P0CA0),
				.a7(P0CB0),
				.a8(P0CC0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00AA2)
);

ninexnine_unit ninexnine_unit_1627(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AA1),
				.a1(P0AB1),
				.a2(P0AC1),
				.a3(P0BA1),
				.a4(P0BB1),
				.a5(P0BC1),
				.a6(P0CA1),
				.a7(P0CB1),
				.a8(P0CC1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01AA2)
);

ninexnine_unit ninexnine_unit_1628(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AA2),
				.a1(P0AB2),
				.a2(P0AC2),
				.a3(P0BA2),
				.a4(P0BB2),
				.a5(P0BC2),
				.a6(P0CA2),
				.a7(P0CB2),
				.a8(P0CC2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02AA2)
);

assign C0AA2=c00AA2+c01AA2+c02AA2;
assign A0AA2=(C0AA2>=0)?1:0;

ninexnine_unit ninexnine_unit_1629(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AB0),
				.a1(P0AC0),
				.a2(P0AD0),
				.a3(P0BB0),
				.a4(P0BC0),
				.a5(P0BD0),
				.a6(P0CB0),
				.a7(P0CC0),
				.a8(P0CD0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00AB2)
);

ninexnine_unit ninexnine_unit_1630(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AB1),
				.a1(P0AC1),
				.a2(P0AD1),
				.a3(P0BB1),
				.a4(P0BC1),
				.a5(P0BD1),
				.a6(P0CB1),
				.a7(P0CC1),
				.a8(P0CD1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01AB2)
);

ninexnine_unit ninexnine_unit_1631(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AB2),
				.a1(P0AC2),
				.a2(P0AD2),
				.a3(P0BB2),
				.a4(P0BC2),
				.a5(P0BD2),
				.a6(P0CB2),
				.a7(P0CC2),
				.a8(P0CD2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02AB2)
);

assign C0AB2=c00AB2+c01AB2+c02AB2;
assign A0AB2=(C0AB2>=0)?1:0;

ninexnine_unit ninexnine_unit_1632(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AC0),
				.a1(P0AD0),
				.a2(P0AE0),
				.a3(P0BC0),
				.a4(P0BD0),
				.a5(P0BE0),
				.a6(P0CC0),
				.a7(P0CD0),
				.a8(P0CE0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00AC2)
);

ninexnine_unit ninexnine_unit_1633(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AC1),
				.a1(P0AD1),
				.a2(P0AE1),
				.a3(P0BC1),
				.a4(P0BD1),
				.a5(P0BE1),
				.a6(P0CC1),
				.a7(P0CD1),
				.a8(P0CE1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01AC2)
);

ninexnine_unit ninexnine_unit_1634(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AC2),
				.a1(P0AD2),
				.a2(P0AE2),
				.a3(P0BC2),
				.a4(P0BD2),
				.a5(P0BE2),
				.a6(P0CC2),
				.a7(P0CD2),
				.a8(P0CE2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02AC2)
);

assign C0AC2=c00AC2+c01AC2+c02AC2;
assign A0AC2=(C0AC2>=0)?1:0;

ninexnine_unit ninexnine_unit_1635(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AD0),
				.a1(P0AE0),
				.a2(P0AF0),
				.a3(P0BD0),
				.a4(P0BE0),
				.a5(P0BF0),
				.a6(P0CD0),
				.a7(P0CE0),
				.a8(P0CF0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00AD2)
);

ninexnine_unit ninexnine_unit_1636(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AD1),
				.a1(P0AE1),
				.a2(P0AF1),
				.a3(P0BD1),
				.a4(P0BE1),
				.a5(P0BF1),
				.a6(P0CD1),
				.a7(P0CE1),
				.a8(P0CF1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01AD2)
);

ninexnine_unit ninexnine_unit_1637(
				.clk(clk),
				.rstn(rstn),
				.a0(P0AD2),
				.a1(P0AE2),
				.a2(P0AF2),
				.a3(P0BD2),
				.a4(P0BE2),
				.a5(P0BF2),
				.a6(P0CD2),
				.a7(P0CE2),
				.a8(P0CF2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02AD2)
);

assign C0AD2=c00AD2+c01AD2+c02AD2;
assign A0AD2=(C0AD2>=0)?1:0;

ninexnine_unit ninexnine_unit_1638(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B00),
				.a1(P0B10),
				.a2(P0B20),
				.a3(P0C00),
				.a4(P0C10),
				.a5(P0C20),
				.a6(P0D00),
				.a7(P0D10),
				.a8(P0D20),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00B02)
);

ninexnine_unit ninexnine_unit_1639(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B01),
				.a1(P0B11),
				.a2(P0B21),
				.a3(P0C01),
				.a4(P0C11),
				.a5(P0C21),
				.a6(P0D01),
				.a7(P0D11),
				.a8(P0D21),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01B02)
);

ninexnine_unit ninexnine_unit_1640(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B02),
				.a1(P0B12),
				.a2(P0B22),
				.a3(P0C02),
				.a4(P0C12),
				.a5(P0C22),
				.a6(P0D02),
				.a7(P0D12),
				.a8(P0D22),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02B02)
);

assign C0B02=c00B02+c01B02+c02B02;
assign A0B02=(C0B02>=0)?1:0;

ninexnine_unit ninexnine_unit_1641(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B10),
				.a1(P0B20),
				.a2(P0B30),
				.a3(P0C10),
				.a4(P0C20),
				.a5(P0C30),
				.a6(P0D10),
				.a7(P0D20),
				.a8(P0D30),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00B12)
);

ninexnine_unit ninexnine_unit_1642(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B11),
				.a1(P0B21),
				.a2(P0B31),
				.a3(P0C11),
				.a4(P0C21),
				.a5(P0C31),
				.a6(P0D11),
				.a7(P0D21),
				.a8(P0D31),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01B12)
);

ninexnine_unit ninexnine_unit_1643(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B12),
				.a1(P0B22),
				.a2(P0B32),
				.a3(P0C12),
				.a4(P0C22),
				.a5(P0C32),
				.a6(P0D12),
				.a7(P0D22),
				.a8(P0D32),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02B12)
);

assign C0B12=c00B12+c01B12+c02B12;
assign A0B12=(C0B12>=0)?1:0;

ninexnine_unit ninexnine_unit_1644(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B20),
				.a1(P0B30),
				.a2(P0B40),
				.a3(P0C20),
				.a4(P0C30),
				.a5(P0C40),
				.a6(P0D20),
				.a7(P0D30),
				.a8(P0D40),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00B22)
);

ninexnine_unit ninexnine_unit_1645(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B21),
				.a1(P0B31),
				.a2(P0B41),
				.a3(P0C21),
				.a4(P0C31),
				.a5(P0C41),
				.a6(P0D21),
				.a7(P0D31),
				.a8(P0D41),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01B22)
);

ninexnine_unit ninexnine_unit_1646(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B22),
				.a1(P0B32),
				.a2(P0B42),
				.a3(P0C22),
				.a4(P0C32),
				.a5(P0C42),
				.a6(P0D22),
				.a7(P0D32),
				.a8(P0D42),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02B22)
);

assign C0B22=c00B22+c01B22+c02B22;
assign A0B22=(C0B22>=0)?1:0;

ninexnine_unit ninexnine_unit_1647(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B30),
				.a1(P0B40),
				.a2(P0B50),
				.a3(P0C30),
				.a4(P0C40),
				.a5(P0C50),
				.a6(P0D30),
				.a7(P0D40),
				.a8(P0D50),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00B32)
);

ninexnine_unit ninexnine_unit_1648(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B31),
				.a1(P0B41),
				.a2(P0B51),
				.a3(P0C31),
				.a4(P0C41),
				.a5(P0C51),
				.a6(P0D31),
				.a7(P0D41),
				.a8(P0D51),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01B32)
);

ninexnine_unit ninexnine_unit_1649(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B32),
				.a1(P0B42),
				.a2(P0B52),
				.a3(P0C32),
				.a4(P0C42),
				.a5(P0C52),
				.a6(P0D32),
				.a7(P0D42),
				.a8(P0D52),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02B32)
);

assign C0B32=c00B32+c01B32+c02B32;
assign A0B32=(C0B32>=0)?1:0;

ninexnine_unit ninexnine_unit_1650(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B40),
				.a1(P0B50),
				.a2(P0B60),
				.a3(P0C40),
				.a4(P0C50),
				.a5(P0C60),
				.a6(P0D40),
				.a7(P0D50),
				.a8(P0D60),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00B42)
);

ninexnine_unit ninexnine_unit_1651(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B41),
				.a1(P0B51),
				.a2(P0B61),
				.a3(P0C41),
				.a4(P0C51),
				.a5(P0C61),
				.a6(P0D41),
				.a7(P0D51),
				.a8(P0D61),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01B42)
);

ninexnine_unit ninexnine_unit_1652(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B42),
				.a1(P0B52),
				.a2(P0B62),
				.a3(P0C42),
				.a4(P0C52),
				.a5(P0C62),
				.a6(P0D42),
				.a7(P0D52),
				.a8(P0D62),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02B42)
);

assign C0B42=c00B42+c01B42+c02B42;
assign A0B42=(C0B42>=0)?1:0;

ninexnine_unit ninexnine_unit_1653(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B50),
				.a1(P0B60),
				.a2(P0B70),
				.a3(P0C50),
				.a4(P0C60),
				.a5(P0C70),
				.a6(P0D50),
				.a7(P0D60),
				.a8(P0D70),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00B52)
);

ninexnine_unit ninexnine_unit_1654(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B51),
				.a1(P0B61),
				.a2(P0B71),
				.a3(P0C51),
				.a4(P0C61),
				.a5(P0C71),
				.a6(P0D51),
				.a7(P0D61),
				.a8(P0D71),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01B52)
);

ninexnine_unit ninexnine_unit_1655(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B52),
				.a1(P0B62),
				.a2(P0B72),
				.a3(P0C52),
				.a4(P0C62),
				.a5(P0C72),
				.a6(P0D52),
				.a7(P0D62),
				.a8(P0D72),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02B52)
);

assign C0B52=c00B52+c01B52+c02B52;
assign A0B52=(C0B52>=0)?1:0;

ninexnine_unit ninexnine_unit_1656(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B60),
				.a1(P0B70),
				.a2(P0B80),
				.a3(P0C60),
				.a4(P0C70),
				.a5(P0C80),
				.a6(P0D60),
				.a7(P0D70),
				.a8(P0D80),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00B62)
);

ninexnine_unit ninexnine_unit_1657(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B61),
				.a1(P0B71),
				.a2(P0B81),
				.a3(P0C61),
				.a4(P0C71),
				.a5(P0C81),
				.a6(P0D61),
				.a7(P0D71),
				.a8(P0D81),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01B62)
);

ninexnine_unit ninexnine_unit_1658(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B62),
				.a1(P0B72),
				.a2(P0B82),
				.a3(P0C62),
				.a4(P0C72),
				.a5(P0C82),
				.a6(P0D62),
				.a7(P0D72),
				.a8(P0D82),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02B62)
);

assign C0B62=c00B62+c01B62+c02B62;
assign A0B62=(C0B62>=0)?1:0;

ninexnine_unit ninexnine_unit_1659(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B70),
				.a1(P0B80),
				.a2(P0B90),
				.a3(P0C70),
				.a4(P0C80),
				.a5(P0C90),
				.a6(P0D70),
				.a7(P0D80),
				.a8(P0D90),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00B72)
);

ninexnine_unit ninexnine_unit_1660(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B71),
				.a1(P0B81),
				.a2(P0B91),
				.a3(P0C71),
				.a4(P0C81),
				.a5(P0C91),
				.a6(P0D71),
				.a7(P0D81),
				.a8(P0D91),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01B72)
);

ninexnine_unit ninexnine_unit_1661(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B72),
				.a1(P0B82),
				.a2(P0B92),
				.a3(P0C72),
				.a4(P0C82),
				.a5(P0C92),
				.a6(P0D72),
				.a7(P0D82),
				.a8(P0D92),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02B72)
);

assign C0B72=c00B72+c01B72+c02B72;
assign A0B72=(C0B72>=0)?1:0;

ninexnine_unit ninexnine_unit_1662(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B80),
				.a1(P0B90),
				.a2(P0BA0),
				.a3(P0C80),
				.a4(P0C90),
				.a5(P0CA0),
				.a6(P0D80),
				.a7(P0D90),
				.a8(P0DA0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00B82)
);

ninexnine_unit ninexnine_unit_1663(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B81),
				.a1(P0B91),
				.a2(P0BA1),
				.a3(P0C81),
				.a4(P0C91),
				.a5(P0CA1),
				.a6(P0D81),
				.a7(P0D91),
				.a8(P0DA1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01B82)
);

ninexnine_unit ninexnine_unit_1664(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B82),
				.a1(P0B92),
				.a2(P0BA2),
				.a3(P0C82),
				.a4(P0C92),
				.a5(P0CA2),
				.a6(P0D82),
				.a7(P0D92),
				.a8(P0DA2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02B82)
);

assign C0B82=c00B82+c01B82+c02B82;
assign A0B82=(C0B82>=0)?1:0;

ninexnine_unit ninexnine_unit_1665(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B90),
				.a1(P0BA0),
				.a2(P0BB0),
				.a3(P0C90),
				.a4(P0CA0),
				.a5(P0CB0),
				.a6(P0D90),
				.a7(P0DA0),
				.a8(P0DB0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00B92)
);

ninexnine_unit ninexnine_unit_1666(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B91),
				.a1(P0BA1),
				.a2(P0BB1),
				.a3(P0C91),
				.a4(P0CA1),
				.a5(P0CB1),
				.a6(P0D91),
				.a7(P0DA1),
				.a8(P0DB1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01B92)
);

ninexnine_unit ninexnine_unit_1667(
				.clk(clk),
				.rstn(rstn),
				.a0(P0B92),
				.a1(P0BA2),
				.a2(P0BB2),
				.a3(P0C92),
				.a4(P0CA2),
				.a5(P0CB2),
				.a6(P0D92),
				.a7(P0DA2),
				.a8(P0DB2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02B92)
);

assign C0B92=c00B92+c01B92+c02B92;
assign A0B92=(C0B92>=0)?1:0;

ninexnine_unit ninexnine_unit_1668(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BA0),
				.a1(P0BB0),
				.a2(P0BC0),
				.a3(P0CA0),
				.a4(P0CB0),
				.a5(P0CC0),
				.a6(P0DA0),
				.a7(P0DB0),
				.a8(P0DC0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00BA2)
);

ninexnine_unit ninexnine_unit_1669(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BA1),
				.a1(P0BB1),
				.a2(P0BC1),
				.a3(P0CA1),
				.a4(P0CB1),
				.a5(P0CC1),
				.a6(P0DA1),
				.a7(P0DB1),
				.a8(P0DC1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01BA2)
);

ninexnine_unit ninexnine_unit_1670(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BA2),
				.a1(P0BB2),
				.a2(P0BC2),
				.a3(P0CA2),
				.a4(P0CB2),
				.a5(P0CC2),
				.a6(P0DA2),
				.a7(P0DB2),
				.a8(P0DC2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02BA2)
);

assign C0BA2=c00BA2+c01BA2+c02BA2;
assign A0BA2=(C0BA2>=0)?1:0;

ninexnine_unit ninexnine_unit_1671(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BB0),
				.a1(P0BC0),
				.a2(P0BD0),
				.a3(P0CB0),
				.a4(P0CC0),
				.a5(P0CD0),
				.a6(P0DB0),
				.a7(P0DC0),
				.a8(P0DD0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00BB2)
);

ninexnine_unit ninexnine_unit_1672(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BB1),
				.a1(P0BC1),
				.a2(P0BD1),
				.a3(P0CB1),
				.a4(P0CC1),
				.a5(P0CD1),
				.a6(P0DB1),
				.a7(P0DC1),
				.a8(P0DD1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01BB2)
);

ninexnine_unit ninexnine_unit_1673(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BB2),
				.a1(P0BC2),
				.a2(P0BD2),
				.a3(P0CB2),
				.a4(P0CC2),
				.a5(P0CD2),
				.a6(P0DB2),
				.a7(P0DC2),
				.a8(P0DD2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02BB2)
);

assign C0BB2=c00BB2+c01BB2+c02BB2;
assign A0BB2=(C0BB2>=0)?1:0;

ninexnine_unit ninexnine_unit_1674(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BC0),
				.a1(P0BD0),
				.a2(P0BE0),
				.a3(P0CC0),
				.a4(P0CD0),
				.a5(P0CE0),
				.a6(P0DC0),
				.a7(P0DD0),
				.a8(P0DE0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00BC2)
);

ninexnine_unit ninexnine_unit_1675(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BC1),
				.a1(P0BD1),
				.a2(P0BE1),
				.a3(P0CC1),
				.a4(P0CD1),
				.a5(P0CE1),
				.a6(P0DC1),
				.a7(P0DD1),
				.a8(P0DE1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01BC2)
);

ninexnine_unit ninexnine_unit_1676(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BC2),
				.a1(P0BD2),
				.a2(P0BE2),
				.a3(P0CC2),
				.a4(P0CD2),
				.a5(P0CE2),
				.a6(P0DC2),
				.a7(P0DD2),
				.a8(P0DE2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02BC2)
);

assign C0BC2=c00BC2+c01BC2+c02BC2;
assign A0BC2=(C0BC2>=0)?1:0;

ninexnine_unit ninexnine_unit_1677(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BD0),
				.a1(P0BE0),
				.a2(P0BF0),
				.a3(P0CD0),
				.a4(P0CE0),
				.a5(P0CF0),
				.a6(P0DD0),
				.a7(P0DE0),
				.a8(P0DF0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00BD2)
);

ninexnine_unit ninexnine_unit_1678(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BD1),
				.a1(P0BE1),
				.a2(P0BF1),
				.a3(P0CD1),
				.a4(P0CE1),
				.a5(P0CF1),
				.a6(P0DD1),
				.a7(P0DE1),
				.a8(P0DF1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01BD2)
);

ninexnine_unit ninexnine_unit_1679(
				.clk(clk),
				.rstn(rstn),
				.a0(P0BD2),
				.a1(P0BE2),
				.a2(P0BF2),
				.a3(P0CD2),
				.a4(P0CE2),
				.a5(P0CF2),
				.a6(P0DD2),
				.a7(P0DE2),
				.a8(P0DF2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02BD2)
);

assign C0BD2=c00BD2+c01BD2+c02BD2;
assign A0BD2=(C0BD2>=0)?1:0;

ninexnine_unit ninexnine_unit_1680(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C00),
				.a1(P0C10),
				.a2(P0C20),
				.a3(P0D00),
				.a4(P0D10),
				.a5(P0D20),
				.a6(P0E00),
				.a7(P0E10),
				.a8(P0E20),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00C02)
);

ninexnine_unit ninexnine_unit_1681(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C01),
				.a1(P0C11),
				.a2(P0C21),
				.a3(P0D01),
				.a4(P0D11),
				.a5(P0D21),
				.a6(P0E01),
				.a7(P0E11),
				.a8(P0E21),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01C02)
);

ninexnine_unit ninexnine_unit_1682(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C02),
				.a1(P0C12),
				.a2(P0C22),
				.a3(P0D02),
				.a4(P0D12),
				.a5(P0D22),
				.a6(P0E02),
				.a7(P0E12),
				.a8(P0E22),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02C02)
);

assign C0C02=c00C02+c01C02+c02C02;
assign A0C02=(C0C02>=0)?1:0;

ninexnine_unit ninexnine_unit_1683(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C10),
				.a1(P0C20),
				.a2(P0C30),
				.a3(P0D10),
				.a4(P0D20),
				.a5(P0D30),
				.a6(P0E10),
				.a7(P0E20),
				.a8(P0E30),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00C12)
);

ninexnine_unit ninexnine_unit_1684(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C11),
				.a1(P0C21),
				.a2(P0C31),
				.a3(P0D11),
				.a4(P0D21),
				.a5(P0D31),
				.a6(P0E11),
				.a7(P0E21),
				.a8(P0E31),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01C12)
);

ninexnine_unit ninexnine_unit_1685(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C12),
				.a1(P0C22),
				.a2(P0C32),
				.a3(P0D12),
				.a4(P0D22),
				.a5(P0D32),
				.a6(P0E12),
				.a7(P0E22),
				.a8(P0E32),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02C12)
);

assign C0C12=c00C12+c01C12+c02C12;
assign A0C12=(C0C12>=0)?1:0;

ninexnine_unit ninexnine_unit_1686(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C20),
				.a1(P0C30),
				.a2(P0C40),
				.a3(P0D20),
				.a4(P0D30),
				.a5(P0D40),
				.a6(P0E20),
				.a7(P0E30),
				.a8(P0E40),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00C22)
);

ninexnine_unit ninexnine_unit_1687(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C21),
				.a1(P0C31),
				.a2(P0C41),
				.a3(P0D21),
				.a4(P0D31),
				.a5(P0D41),
				.a6(P0E21),
				.a7(P0E31),
				.a8(P0E41),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01C22)
);

ninexnine_unit ninexnine_unit_1688(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C22),
				.a1(P0C32),
				.a2(P0C42),
				.a3(P0D22),
				.a4(P0D32),
				.a5(P0D42),
				.a6(P0E22),
				.a7(P0E32),
				.a8(P0E42),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02C22)
);

assign C0C22=c00C22+c01C22+c02C22;
assign A0C22=(C0C22>=0)?1:0;

ninexnine_unit ninexnine_unit_1689(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C30),
				.a1(P0C40),
				.a2(P0C50),
				.a3(P0D30),
				.a4(P0D40),
				.a5(P0D50),
				.a6(P0E30),
				.a7(P0E40),
				.a8(P0E50),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00C32)
);

ninexnine_unit ninexnine_unit_1690(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C31),
				.a1(P0C41),
				.a2(P0C51),
				.a3(P0D31),
				.a4(P0D41),
				.a5(P0D51),
				.a6(P0E31),
				.a7(P0E41),
				.a8(P0E51),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01C32)
);

ninexnine_unit ninexnine_unit_1691(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C32),
				.a1(P0C42),
				.a2(P0C52),
				.a3(P0D32),
				.a4(P0D42),
				.a5(P0D52),
				.a6(P0E32),
				.a7(P0E42),
				.a8(P0E52),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02C32)
);

assign C0C32=c00C32+c01C32+c02C32;
assign A0C32=(C0C32>=0)?1:0;

ninexnine_unit ninexnine_unit_1692(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C40),
				.a1(P0C50),
				.a2(P0C60),
				.a3(P0D40),
				.a4(P0D50),
				.a5(P0D60),
				.a6(P0E40),
				.a7(P0E50),
				.a8(P0E60),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00C42)
);

ninexnine_unit ninexnine_unit_1693(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C41),
				.a1(P0C51),
				.a2(P0C61),
				.a3(P0D41),
				.a4(P0D51),
				.a5(P0D61),
				.a6(P0E41),
				.a7(P0E51),
				.a8(P0E61),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01C42)
);

ninexnine_unit ninexnine_unit_1694(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C42),
				.a1(P0C52),
				.a2(P0C62),
				.a3(P0D42),
				.a4(P0D52),
				.a5(P0D62),
				.a6(P0E42),
				.a7(P0E52),
				.a8(P0E62),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02C42)
);

assign C0C42=c00C42+c01C42+c02C42;
assign A0C42=(C0C42>=0)?1:0;

ninexnine_unit ninexnine_unit_1695(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C50),
				.a1(P0C60),
				.a2(P0C70),
				.a3(P0D50),
				.a4(P0D60),
				.a5(P0D70),
				.a6(P0E50),
				.a7(P0E60),
				.a8(P0E70),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00C52)
);

ninexnine_unit ninexnine_unit_1696(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C51),
				.a1(P0C61),
				.a2(P0C71),
				.a3(P0D51),
				.a4(P0D61),
				.a5(P0D71),
				.a6(P0E51),
				.a7(P0E61),
				.a8(P0E71),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01C52)
);

ninexnine_unit ninexnine_unit_1697(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C52),
				.a1(P0C62),
				.a2(P0C72),
				.a3(P0D52),
				.a4(P0D62),
				.a5(P0D72),
				.a6(P0E52),
				.a7(P0E62),
				.a8(P0E72),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02C52)
);

assign C0C52=c00C52+c01C52+c02C52;
assign A0C52=(C0C52>=0)?1:0;

ninexnine_unit ninexnine_unit_1698(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C60),
				.a1(P0C70),
				.a2(P0C80),
				.a3(P0D60),
				.a4(P0D70),
				.a5(P0D80),
				.a6(P0E60),
				.a7(P0E70),
				.a8(P0E80),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00C62)
);

ninexnine_unit ninexnine_unit_1699(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C61),
				.a1(P0C71),
				.a2(P0C81),
				.a3(P0D61),
				.a4(P0D71),
				.a5(P0D81),
				.a6(P0E61),
				.a7(P0E71),
				.a8(P0E81),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01C62)
);

ninexnine_unit ninexnine_unit_1700(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C62),
				.a1(P0C72),
				.a2(P0C82),
				.a3(P0D62),
				.a4(P0D72),
				.a5(P0D82),
				.a6(P0E62),
				.a7(P0E72),
				.a8(P0E82),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02C62)
);

assign C0C62=c00C62+c01C62+c02C62;
assign A0C62=(C0C62>=0)?1:0;

ninexnine_unit ninexnine_unit_1701(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C70),
				.a1(P0C80),
				.a2(P0C90),
				.a3(P0D70),
				.a4(P0D80),
				.a5(P0D90),
				.a6(P0E70),
				.a7(P0E80),
				.a8(P0E90),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00C72)
);

ninexnine_unit ninexnine_unit_1702(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C71),
				.a1(P0C81),
				.a2(P0C91),
				.a3(P0D71),
				.a4(P0D81),
				.a5(P0D91),
				.a6(P0E71),
				.a7(P0E81),
				.a8(P0E91),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01C72)
);

ninexnine_unit ninexnine_unit_1703(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C72),
				.a1(P0C82),
				.a2(P0C92),
				.a3(P0D72),
				.a4(P0D82),
				.a5(P0D92),
				.a6(P0E72),
				.a7(P0E82),
				.a8(P0E92),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02C72)
);

assign C0C72=c00C72+c01C72+c02C72;
assign A0C72=(C0C72>=0)?1:0;

ninexnine_unit ninexnine_unit_1704(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C80),
				.a1(P0C90),
				.a2(P0CA0),
				.a3(P0D80),
				.a4(P0D90),
				.a5(P0DA0),
				.a6(P0E80),
				.a7(P0E90),
				.a8(P0EA0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00C82)
);

ninexnine_unit ninexnine_unit_1705(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C81),
				.a1(P0C91),
				.a2(P0CA1),
				.a3(P0D81),
				.a4(P0D91),
				.a5(P0DA1),
				.a6(P0E81),
				.a7(P0E91),
				.a8(P0EA1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01C82)
);

ninexnine_unit ninexnine_unit_1706(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C82),
				.a1(P0C92),
				.a2(P0CA2),
				.a3(P0D82),
				.a4(P0D92),
				.a5(P0DA2),
				.a6(P0E82),
				.a7(P0E92),
				.a8(P0EA2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02C82)
);

assign C0C82=c00C82+c01C82+c02C82;
assign A0C82=(C0C82>=0)?1:0;

ninexnine_unit ninexnine_unit_1707(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C90),
				.a1(P0CA0),
				.a2(P0CB0),
				.a3(P0D90),
				.a4(P0DA0),
				.a5(P0DB0),
				.a6(P0E90),
				.a7(P0EA0),
				.a8(P0EB0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00C92)
);

ninexnine_unit ninexnine_unit_1708(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C91),
				.a1(P0CA1),
				.a2(P0CB1),
				.a3(P0D91),
				.a4(P0DA1),
				.a5(P0DB1),
				.a6(P0E91),
				.a7(P0EA1),
				.a8(P0EB1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01C92)
);

ninexnine_unit ninexnine_unit_1709(
				.clk(clk),
				.rstn(rstn),
				.a0(P0C92),
				.a1(P0CA2),
				.a2(P0CB2),
				.a3(P0D92),
				.a4(P0DA2),
				.a5(P0DB2),
				.a6(P0E92),
				.a7(P0EA2),
				.a8(P0EB2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02C92)
);

assign C0C92=c00C92+c01C92+c02C92;
assign A0C92=(C0C92>=0)?1:0;

ninexnine_unit ninexnine_unit_1710(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CA0),
				.a1(P0CB0),
				.a2(P0CC0),
				.a3(P0DA0),
				.a4(P0DB0),
				.a5(P0DC0),
				.a6(P0EA0),
				.a7(P0EB0),
				.a8(P0EC0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00CA2)
);

ninexnine_unit ninexnine_unit_1711(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CA1),
				.a1(P0CB1),
				.a2(P0CC1),
				.a3(P0DA1),
				.a4(P0DB1),
				.a5(P0DC1),
				.a6(P0EA1),
				.a7(P0EB1),
				.a8(P0EC1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01CA2)
);

ninexnine_unit ninexnine_unit_1712(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CA2),
				.a1(P0CB2),
				.a2(P0CC2),
				.a3(P0DA2),
				.a4(P0DB2),
				.a5(P0DC2),
				.a6(P0EA2),
				.a7(P0EB2),
				.a8(P0EC2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02CA2)
);

assign C0CA2=c00CA2+c01CA2+c02CA2;
assign A0CA2=(C0CA2>=0)?1:0;

ninexnine_unit ninexnine_unit_1713(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CB0),
				.a1(P0CC0),
				.a2(P0CD0),
				.a3(P0DB0),
				.a4(P0DC0),
				.a5(P0DD0),
				.a6(P0EB0),
				.a7(P0EC0),
				.a8(P0ED0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00CB2)
);

ninexnine_unit ninexnine_unit_1714(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CB1),
				.a1(P0CC1),
				.a2(P0CD1),
				.a3(P0DB1),
				.a4(P0DC1),
				.a5(P0DD1),
				.a6(P0EB1),
				.a7(P0EC1),
				.a8(P0ED1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01CB2)
);

ninexnine_unit ninexnine_unit_1715(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CB2),
				.a1(P0CC2),
				.a2(P0CD2),
				.a3(P0DB2),
				.a4(P0DC2),
				.a5(P0DD2),
				.a6(P0EB2),
				.a7(P0EC2),
				.a8(P0ED2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02CB2)
);

assign C0CB2=c00CB2+c01CB2+c02CB2;
assign A0CB2=(C0CB2>=0)?1:0;

ninexnine_unit ninexnine_unit_1716(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CC0),
				.a1(P0CD0),
				.a2(P0CE0),
				.a3(P0DC0),
				.a4(P0DD0),
				.a5(P0DE0),
				.a6(P0EC0),
				.a7(P0ED0),
				.a8(P0EE0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00CC2)
);

ninexnine_unit ninexnine_unit_1717(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CC1),
				.a1(P0CD1),
				.a2(P0CE1),
				.a3(P0DC1),
				.a4(P0DD1),
				.a5(P0DE1),
				.a6(P0EC1),
				.a7(P0ED1),
				.a8(P0EE1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01CC2)
);

ninexnine_unit ninexnine_unit_1718(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CC2),
				.a1(P0CD2),
				.a2(P0CE2),
				.a3(P0DC2),
				.a4(P0DD2),
				.a5(P0DE2),
				.a6(P0EC2),
				.a7(P0ED2),
				.a8(P0EE2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02CC2)
);

assign C0CC2=c00CC2+c01CC2+c02CC2;
assign A0CC2=(C0CC2>=0)?1:0;

ninexnine_unit ninexnine_unit_1719(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CD0),
				.a1(P0CE0),
				.a2(P0CF0),
				.a3(P0DD0),
				.a4(P0DE0),
				.a5(P0DF0),
				.a6(P0ED0),
				.a7(P0EE0),
				.a8(P0EF0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00CD2)
);

ninexnine_unit ninexnine_unit_1720(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CD1),
				.a1(P0CE1),
				.a2(P0CF1),
				.a3(P0DD1),
				.a4(P0DE1),
				.a5(P0DF1),
				.a6(P0ED1),
				.a7(P0EE1),
				.a8(P0EF1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01CD2)
);

ninexnine_unit ninexnine_unit_1721(
				.clk(clk),
				.rstn(rstn),
				.a0(P0CD2),
				.a1(P0CE2),
				.a2(P0CF2),
				.a3(P0DD2),
				.a4(P0DE2),
				.a5(P0DF2),
				.a6(P0ED2),
				.a7(P0EE2),
				.a8(P0EF2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02CD2)
);

assign C0CD2=c00CD2+c01CD2+c02CD2;
assign A0CD2=(C0CD2>=0)?1:0;

ninexnine_unit ninexnine_unit_1722(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D00),
				.a1(P0D10),
				.a2(P0D20),
				.a3(P0E00),
				.a4(P0E10),
				.a5(P0E20),
				.a6(P0F00),
				.a7(P0F10),
				.a8(P0F20),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00D02)
);

ninexnine_unit ninexnine_unit_1723(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D01),
				.a1(P0D11),
				.a2(P0D21),
				.a3(P0E01),
				.a4(P0E11),
				.a5(P0E21),
				.a6(P0F01),
				.a7(P0F11),
				.a8(P0F21),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01D02)
);

ninexnine_unit ninexnine_unit_1724(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D02),
				.a1(P0D12),
				.a2(P0D22),
				.a3(P0E02),
				.a4(P0E12),
				.a5(P0E22),
				.a6(P0F02),
				.a7(P0F12),
				.a8(P0F22),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02D02)
);

assign C0D02=c00D02+c01D02+c02D02;
assign A0D02=(C0D02>=0)?1:0;

ninexnine_unit ninexnine_unit_1725(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D10),
				.a1(P0D20),
				.a2(P0D30),
				.a3(P0E10),
				.a4(P0E20),
				.a5(P0E30),
				.a6(P0F10),
				.a7(P0F20),
				.a8(P0F30),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00D12)
);

ninexnine_unit ninexnine_unit_1726(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D11),
				.a1(P0D21),
				.a2(P0D31),
				.a3(P0E11),
				.a4(P0E21),
				.a5(P0E31),
				.a6(P0F11),
				.a7(P0F21),
				.a8(P0F31),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01D12)
);

ninexnine_unit ninexnine_unit_1727(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D12),
				.a1(P0D22),
				.a2(P0D32),
				.a3(P0E12),
				.a4(P0E22),
				.a5(P0E32),
				.a6(P0F12),
				.a7(P0F22),
				.a8(P0F32),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02D12)
);

assign C0D12=c00D12+c01D12+c02D12;
assign A0D12=(C0D12>=0)?1:0;

ninexnine_unit ninexnine_unit_1728(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D20),
				.a1(P0D30),
				.a2(P0D40),
				.a3(P0E20),
				.a4(P0E30),
				.a5(P0E40),
				.a6(P0F20),
				.a7(P0F30),
				.a8(P0F40),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00D22)
);

ninexnine_unit ninexnine_unit_1729(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D21),
				.a1(P0D31),
				.a2(P0D41),
				.a3(P0E21),
				.a4(P0E31),
				.a5(P0E41),
				.a6(P0F21),
				.a7(P0F31),
				.a8(P0F41),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01D22)
);

ninexnine_unit ninexnine_unit_1730(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D22),
				.a1(P0D32),
				.a2(P0D42),
				.a3(P0E22),
				.a4(P0E32),
				.a5(P0E42),
				.a6(P0F22),
				.a7(P0F32),
				.a8(P0F42),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02D22)
);

assign C0D22=c00D22+c01D22+c02D22;
assign A0D22=(C0D22>=0)?1:0;

ninexnine_unit ninexnine_unit_1731(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D30),
				.a1(P0D40),
				.a2(P0D50),
				.a3(P0E30),
				.a4(P0E40),
				.a5(P0E50),
				.a6(P0F30),
				.a7(P0F40),
				.a8(P0F50),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00D32)
);

ninexnine_unit ninexnine_unit_1732(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D31),
				.a1(P0D41),
				.a2(P0D51),
				.a3(P0E31),
				.a4(P0E41),
				.a5(P0E51),
				.a6(P0F31),
				.a7(P0F41),
				.a8(P0F51),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01D32)
);

ninexnine_unit ninexnine_unit_1733(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D32),
				.a1(P0D42),
				.a2(P0D52),
				.a3(P0E32),
				.a4(P0E42),
				.a5(P0E52),
				.a6(P0F32),
				.a7(P0F42),
				.a8(P0F52),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02D32)
);

assign C0D32=c00D32+c01D32+c02D32;
assign A0D32=(C0D32>=0)?1:0;

ninexnine_unit ninexnine_unit_1734(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D40),
				.a1(P0D50),
				.a2(P0D60),
				.a3(P0E40),
				.a4(P0E50),
				.a5(P0E60),
				.a6(P0F40),
				.a7(P0F50),
				.a8(P0F60),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00D42)
);

ninexnine_unit ninexnine_unit_1735(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D41),
				.a1(P0D51),
				.a2(P0D61),
				.a3(P0E41),
				.a4(P0E51),
				.a5(P0E61),
				.a6(P0F41),
				.a7(P0F51),
				.a8(P0F61),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01D42)
);

ninexnine_unit ninexnine_unit_1736(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D42),
				.a1(P0D52),
				.a2(P0D62),
				.a3(P0E42),
				.a4(P0E52),
				.a5(P0E62),
				.a6(P0F42),
				.a7(P0F52),
				.a8(P0F62),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02D42)
);

assign C0D42=c00D42+c01D42+c02D42;
assign A0D42=(C0D42>=0)?1:0;

ninexnine_unit ninexnine_unit_1737(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D50),
				.a1(P0D60),
				.a2(P0D70),
				.a3(P0E50),
				.a4(P0E60),
				.a5(P0E70),
				.a6(P0F50),
				.a7(P0F60),
				.a8(P0F70),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00D52)
);

ninexnine_unit ninexnine_unit_1738(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D51),
				.a1(P0D61),
				.a2(P0D71),
				.a3(P0E51),
				.a4(P0E61),
				.a5(P0E71),
				.a6(P0F51),
				.a7(P0F61),
				.a8(P0F71),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01D52)
);

ninexnine_unit ninexnine_unit_1739(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D52),
				.a1(P0D62),
				.a2(P0D72),
				.a3(P0E52),
				.a4(P0E62),
				.a5(P0E72),
				.a6(P0F52),
				.a7(P0F62),
				.a8(P0F72),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02D52)
);

assign C0D52=c00D52+c01D52+c02D52;
assign A0D52=(C0D52>=0)?1:0;

ninexnine_unit ninexnine_unit_1740(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D60),
				.a1(P0D70),
				.a2(P0D80),
				.a3(P0E60),
				.a4(P0E70),
				.a5(P0E80),
				.a6(P0F60),
				.a7(P0F70),
				.a8(P0F80),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00D62)
);

ninexnine_unit ninexnine_unit_1741(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D61),
				.a1(P0D71),
				.a2(P0D81),
				.a3(P0E61),
				.a4(P0E71),
				.a5(P0E81),
				.a6(P0F61),
				.a7(P0F71),
				.a8(P0F81),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01D62)
);

ninexnine_unit ninexnine_unit_1742(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D62),
				.a1(P0D72),
				.a2(P0D82),
				.a3(P0E62),
				.a4(P0E72),
				.a5(P0E82),
				.a6(P0F62),
				.a7(P0F72),
				.a8(P0F82),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02D62)
);

assign C0D62=c00D62+c01D62+c02D62;
assign A0D62=(C0D62>=0)?1:0;

ninexnine_unit ninexnine_unit_1743(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D70),
				.a1(P0D80),
				.a2(P0D90),
				.a3(P0E70),
				.a4(P0E80),
				.a5(P0E90),
				.a6(P0F70),
				.a7(P0F80),
				.a8(P0F90),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00D72)
);

ninexnine_unit ninexnine_unit_1744(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D71),
				.a1(P0D81),
				.a2(P0D91),
				.a3(P0E71),
				.a4(P0E81),
				.a5(P0E91),
				.a6(P0F71),
				.a7(P0F81),
				.a8(P0F91),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01D72)
);

ninexnine_unit ninexnine_unit_1745(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D72),
				.a1(P0D82),
				.a2(P0D92),
				.a3(P0E72),
				.a4(P0E82),
				.a5(P0E92),
				.a6(P0F72),
				.a7(P0F82),
				.a8(P0F92),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02D72)
);

assign C0D72=c00D72+c01D72+c02D72;
assign A0D72=(C0D72>=0)?1:0;

ninexnine_unit ninexnine_unit_1746(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D80),
				.a1(P0D90),
				.a2(P0DA0),
				.a3(P0E80),
				.a4(P0E90),
				.a5(P0EA0),
				.a6(P0F80),
				.a7(P0F90),
				.a8(P0FA0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00D82)
);

ninexnine_unit ninexnine_unit_1747(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D81),
				.a1(P0D91),
				.a2(P0DA1),
				.a3(P0E81),
				.a4(P0E91),
				.a5(P0EA1),
				.a6(P0F81),
				.a7(P0F91),
				.a8(P0FA1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01D82)
);

ninexnine_unit ninexnine_unit_1748(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D82),
				.a1(P0D92),
				.a2(P0DA2),
				.a3(P0E82),
				.a4(P0E92),
				.a5(P0EA2),
				.a6(P0F82),
				.a7(P0F92),
				.a8(P0FA2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02D82)
);

assign C0D82=c00D82+c01D82+c02D82;
assign A0D82=(C0D82>=0)?1:0;

ninexnine_unit ninexnine_unit_1749(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D90),
				.a1(P0DA0),
				.a2(P0DB0),
				.a3(P0E90),
				.a4(P0EA0),
				.a5(P0EB0),
				.a6(P0F90),
				.a7(P0FA0),
				.a8(P0FB0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00D92)
);

ninexnine_unit ninexnine_unit_1750(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D91),
				.a1(P0DA1),
				.a2(P0DB1),
				.a3(P0E91),
				.a4(P0EA1),
				.a5(P0EB1),
				.a6(P0F91),
				.a7(P0FA1),
				.a8(P0FB1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01D92)
);

ninexnine_unit ninexnine_unit_1751(
				.clk(clk),
				.rstn(rstn),
				.a0(P0D92),
				.a1(P0DA2),
				.a2(P0DB2),
				.a3(P0E92),
				.a4(P0EA2),
				.a5(P0EB2),
				.a6(P0F92),
				.a7(P0FA2),
				.a8(P0FB2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02D92)
);

assign C0D92=c00D92+c01D92+c02D92;
assign A0D92=(C0D92>=0)?1:0;

ninexnine_unit ninexnine_unit_1752(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DA0),
				.a1(P0DB0),
				.a2(P0DC0),
				.a3(P0EA0),
				.a4(P0EB0),
				.a5(P0EC0),
				.a6(P0FA0),
				.a7(P0FB0),
				.a8(P0FC0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00DA2)
);

ninexnine_unit ninexnine_unit_1753(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DA1),
				.a1(P0DB1),
				.a2(P0DC1),
				.a3(P0EA1),
				.a4(P0EB1),
				.a5(P0EC1),
				.a6(P0FA1),
				.a7(P0FB1),
				.a8(P0FC1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01DA2)
);

ninexnine_unit ninexnine_unit_1754(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DA2),
				.a1(P0DB2),
				.a2(P0DC2),
				.a3(P0EA2),
				.a4(P0EB2),
				.a5(P0EC2),
				.a6(P0FA2),
				.a7(P0FB2),
				.a8(P0FC2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02DA2)
);

assign C0DA2=c00DA2+c01DA2+c02DA2;
assign A0DA2=(C0DA2>=0)?1:0;

ninexnine_unit ninexnine_unit_1755(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DB0),
				.a1(P0DC0),
				.a2(P0DD0),
				.a3(P0EB0),
				.a4(P0EC0),
				.a5(P0ED0),
				.a6(P0FB0),
				.a7(P0FC0),
				.a8(P0FD0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00DB2)
);

ninexnine_unit ninexnine_unit_1756(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DB1),
				.a1(P0DC1),
				.a2(P0DD1),
				.a3(P0EB1),
				.a4(P0EC1),
				.a5(P0ED1),
				.a6(P0FB1),
				.a7(P0FC1),
				.a8(P0FD1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01DB2)
);

ninexnine_unit ninexnine_unit_1757(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DB2),
				.a1(P0DC2),
				.a2(P0DD2),
				.a3(P0EB2),
				.a4(P0EC2),
				.a5(P0ED2),
				.a6(P0FB2),
				.a7(P0FC2),
				.a8(P0FD2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02DB2)
);

assign C0DB2=c00DB2+c01DB2+c02DB2;
assign A0DB2=(C0DB2>=0)?1:0;

ninexnine_unit ninexnine_unit_1758(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DC0),
				.a1(P0DD0),
				.a2(P0DE0),
				.a3(P0EC0),
				.a4(P0ED0),
				.a5(P0EE0),
				.a6(P0FC0),
				.a7(P0FD0),
				.a8(P0FE0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00DC2)
);

ninexnine_unit ninexnine_unit_1759(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DC1),
				.a1(P0DD1),
				.a2(P0DE1),
				.a3(P0EC1),
				.a4(P0ED1),
				.a5(P0EE1),
				.a6(P0FC1),
				.a7(P0FD1),
				.a8(P0FE1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01DC2)
);

ninexnine_unit ninexnine_unit_1760(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DC2),
				.a1(P0DD2),
				.a2(P0DE2),
				.a3(P0EC2),
				.a4(P0ED2),
				.a5(P0EE2),
				.a6(P0FC2),
				.a7(P0FD2),
				.a8(P0FE2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02DC2)
);

assign C0DC2=c00DC2+c01DC2+c02DC2;
assign A0DC2=(C0DC2>=0)?1:0;

ninexnine_unit ninexnine_unit_1761(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DD0),
				.a1(P0DE0),
				.a2(P0DF0),
				.a3(P0ED0),
				.a4(P0EE0),
				.a5(P0EF0),
				.a6(P0FD0),
				.a7(P0FE0),
				.a8(P0FF0),
				.b0(W02000),
				.b1(W02010),
				.b2(W02020),
				.b3(W02100),
				.b4(W02110),
				.b5(W02120),
				.b6(W02200),
				.b7(W02210),
				.b8(W02220),
				.c(c00DD2)
);

ninexnine_unit ninexnine_unit_1762(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DD1),
				.a1(P0DE1),
				.a2(P0DF1),
				.a3(P0ED1),
				.a4(P0EE1),
				.a5(P0EF1),
				.a6(P0FD1),
				.a7(P0FE1),
				.a8(P0FF1),
				.b0(W02001),
				.b1(W02011),
				.b2(W02021),
				.b3(W02101),
				.b4(W02111),
				.b5(W02121),
				.b6(W02201),
				.b7(W02211),
				.b8(W02221),
				.c(c01DD2)
);

ninexnine_unit ninexnine_unit_1763(
				.clk(clk),
				.rstn(rstn),
				.a0(P0DD2),
				.a1(P0DE2),
				.a2(P0DF2),
				.a3(P0ED2),
				.a4(P0EE2),
				.a5(P0EF2),
				.a6(P0FD2),
				.a7(P0FE2),
				.a8(P0FF2),
				.b0(W02002),
				.b1(W02012),
				.b2(W02022),
				.b3(W02102),
				.b4(W02112),
				.b5(W02122),
				.b6(W02202),
				.b7(W02212),
				.b8(W02222),
				.c(c02DD2)
);

assign C0DD2=c00DD2+c01DD2+c02DD2;
assign A0DD2=(C0DD2>=0)?1:0;

maxpool maxpool_0(
				.clk(clk),
				.rstn(rstn),
				.a0(A0000),
				.a1(A0010),
				.a2(A0100),
				.a3(A0110),
				.p(P1000)
);

maxpool maxpool_1(
				.clk(clk),
				.rstn(rstn),
				.a0(A0020),
				.a1(A0030),
				.a2(A0120),
				.a3(A0130),
				.p(P1010)
);

maxpool maxpool_2(
				.clk(clk),
				.rstn(rstn),
				.a0(A0040),
				.a1(A0050),
				.a2(A0140),
				.a3(A0150),
				.p(P1020)
);

maxpool maxpool_3(
				.clk(clk),
				.rstn(rstn),
				.a0(A0060),
				.a1(A0070),
				.a2(A0160),
				.a3(A0170),
				.p(P1030)
);

maxpool maxpool_4(
				.clk(clk),
				.rstn(rstn),
				.a0(A0080),
				.a1(A0090),
				.a2(A0180),
				.a3(A0190),
				.p(P1040)
);

maxpool maxpool_5(
				.clk(clk),
				.rstn(rstn),
				.a0(A00A0),
				.a1(A00B0),
				.a2(A01A0),
				.a3(A01B0),
				.p(P1050)
);

maxpool maxpool_6(
				.clk(clk),
				.rstn(rstn),
				.a0(A00C0),
				.a1(A00D0),
				.a2(A01C0),
				.a3(A01D0),
				.p(P1060)
);

maxpool maxpool_7(
				.clk(clk),
				.rstn(rstn),
				.a0(A0200),
				.a1(A0210),
				.a2(A0300),
				.a3(A0310),
				.p(P1100)
);

maxpool maxpool_8(
				.clk(clk),
				.rstn(rstn),
				.a0(A0220),
				.a1(A0230),
				.a2(A0320),
				.a3(A0330),
				.p(P1110)
);

maxpool maxpool_9(
				.clk(clk),
				.rstn(rstn),
				.a0(A0240),
				.a1(A0250),
				.a2(A0340),
				.a3(A0350),
				.p(P1120)
);

maxpool maxpool_10(
				.clk(clk),
				.rstn(rstn),
				.a0(A0260),
				.a1(A0270),
				.a2(A0360),
				.a3(A0370),
				.p(P1130)
);

maxpool maxpool_11(
				.clk(clk),
				.rstn(rstn),
				.a0(A0280),
				.a1(A0290),
				.a2(A0380),
				.a3(A0390),
				.p(P1140)
);

maxpool maxpool_12(
				.clk(clk),
				.rstn(rstn),
				.a0(A02A0),
				.a1(A02B0),
				.a2(A03A0),
				.a3(A03B0),
				.p(P1150)
);

maxpool maxpool_13(
				.clk(clk),
				.rstn(rstn),
				.a0(A02C0),
				.a1(A02D0),
				.a2(A03C0),
				.a3(A03D0),
				.p(P1160)
);

maxpool maxpool_14(
				.clk(clk),
				.rstn(rstn),
				.a0(A0400),
				.a1(A0410),
				.a2(A0500),
				.a3(A0510),
				.p(P1200)
);

maxpool maxpool_15(
				.clk(clk),
				.rstn(rstn),
				.a0(A0420),
				.a1(A0430),
				.a2(A0520),
				.a3(A0530),
				.p(P1210)
);

maxpool maxpool_16(
				.clk(clk),
				.rstn(rstn),
				.a0(A0440),
				.a1(A0450),
				.a2(A0540),
				.a3(A0550),
				.p(P1220)
);

maxpool maxpool_17(
				.clk(clk),
				.rstn(rstn),
				.a0(A0460),
				.a1(A0470),
				.a2(A0560),
				.a3(A0570),
				.p(P1230)
);

maxpool maxpool_18(
				.clk(clk),
				.rstn(rstn),
				.a0(A0480),
				.a1(A0490),
				.a2(A0580),
				.a3(A0590),
				.p(P1240)
);

maxpool maxpool_19(
				.clk(clk),
				.rstn(rstn),
				.a0(A04A0),
				.a1(A04B0),
				.a2(A05A0),
				.a3(A05B0),
				.p(P1250)
);

maxpool maxpool_20(
				.clk(clk),
				.rstn(rstn),
				.a0(A04C0),
				.a1(A04D0),
				.a2(A05C0),
				.a3(A05D0),
				.p(P1260)
);

maxpool maxpool_21(
				.clk(clk),
				.rstn(rstn),
				.a0(A0600),
				.a1(A0610),
				.a2(A0700),
				.a3(A0710),
				.p(P1300)
);

maxpool maxpool_22(
				.clk(clk),
				.rstn(rstn),
				.a0(A0620),
				.a1(A0630),
				.a2(A0720),
				.a3(A0730),
				.p(P1310)
);

maxpool maxpool_23(
				.clk(clk),
				.rstn(rstn),
				.a0(A0640),
				.a1(A0650),
				.a2(A0740),
				.a3(A0750),
				.p(P1320)
);

maxpool maxpool_24(
				.clk(clk),
				.rstn(rstn),
				.a0(A0660),
				.a1(A0670),
				.a2(A0760),
				.a3(A0770),
				.p(P1330)
);

maxpool maxpool_25(
				.clk(clk),
				.rstn(rstn),
				.a0(A0680),
				.a1(A0690),
				.a2(A0780),
				.a3(A0790),
				.p(P1340)
);

maxpool maxpool_26(
				.clk(clk),
				.rstn(rstn),
				.a0(A06A0),
				.a1(A06B0),
				.a2(A07A0),
				.a3(A07B0),
				.p(P1350)
);

maxpool maxpool_27(
				.clk(clk),
				.rstn(rstn),
				.a0(A06C0),
				.a1(A06D0),
				.a2(A07C0),
				.a3(A07D0),
				.p(P1360)
);

maxpool maxpool_28(
				.clk(clk),
				.rstn(rstn),
				.a0(A0800),
				.a1(A0810),
				.a2(A0900),
				.a3(A0910),
				.p(P1400)
);

maxpool maxpool_29(
				.clk(clk),
				.rstn(rstn),
				.a0(A0820),
				.a1(A0830),
				.a2(A0920),
				.a3(A0930),
				.p(P1410)
);

maxpool maxpool_30(
				.clk(clk),
				.rstn(rstn),
				.a0(A0840),
				.a1(A0850),
				.a2(A0940),
				.a3(A0950),
				.p(P1420)
);

maxpool maxpool_31(
				.clk(clk),
				.rstn(rstn),
				.a0(A0860),
				.a1(A0870),
				.a2(A0960),
				.a3(A0970),
				.p(P1430)
);

maxpool maxpool_32(
				.clk(clk),
				.rstn(rstn),
				.a0(A0880),
				.a1(A0890),
				.a2(A0980),
				.a3(A0990),
				.p(P1440)
);

maxpool maxpool_33(
				.clk(clk),
				.rstn(rstn),
				.a0(A08A0),
				.a1(A08B0),
				.a2(A09A0),
				.a3(A09B0),
				.p(P1450)
);

maxpool maxpool_34(
				.clk(clk),
				.rstn(rstn),
				.a0(A08C0),
				.a1(A08D0),
				.a2(A09C0),
				.a3(A09D0),
				.p(P1460)
);

maxpool maxpool_35(
				.clk(clk),
				.rstn(rstn),
				.a0(A0A00),
				.a1(A0A10),
				.a2(A0B00),
				.a3(A0B10),
				.p(P1500)
);

maxpool maxpool_36(
				.clk(clk),
				.rstn(rstn),
				.a0(A0A20),
				.a1(A0A30),
				.a2(A0B20),
				.a3(A0B30),
				.p(P1510)
);

maxpool maxpool_37(
				.clk(clk),
				.rstn(rstn),
				.a0(A0A40),
				.a1(A0A50),
				.a2(A0B40),
				.a3(A0B50),
				.p(P1520)
);

maxpool maxpool_38(
				.clk(clk),
				.rstn(rstn),
				.a0(A0A60),
				.a1(A0A70),
				.a2(A0B60),
				.a3(A0B70),
				.p(P1530)
);

maxpool maxpool_39(
				.clk(clk),
				.rstn(rstn),
				.a0(A0A80),
				.a1(A0A90),
				.a2(A0B80),
				.a3(A0B90),
				.p(P1540)
);

maxpool maxpool_40(
				.clk(clk),
				.rstn(rstn),
				.a0(A0AA0),
				.a1(A0AB0),
				.a2(A0BA0),
				.a3(A0BB0),
				.p(P1550)
);

maxpool maxpool_41(
				.clk(clk),
				.rstn(rstn),
				.a0(A0AC0),
				.a1(A0AD0),
				.a2(A0BC0),
				.a3(A0BD0),
				.p(P1560)
);

maxpool maxpool_42(
				.clk(clk),
				.rstn(rstn),
				.a0(A0C00),
				.a1(A0C10),
				.a2(A0D00),
				.a3(A0D10),
				.p(P1600)
);

maxpool maxpool_43(
				.clk(clk),
				.rstn(rstn),
				.a0(A0C20),
				.a1(A0C30),
				.a2(A0D20),
				.a3(A0D30),
				.p(P1610)
);

maxpool maxpool_44(
				.clk(clk),
				.rstn(rstn),
				.a0(A0C40),
				.a1(A0C50),
				.a2(A0D40),
				.a3(A0D50),
				.p(P1620)
);

maxpool maxpool_45(
				.clk(clk),
				.rstn(rstn),
				.a0(A0C60),
				.a1(A0C70),
				.a2(A0D60),
				.a3(A0D70),
				.p(P1630)
);

maxpool maxpool_46(
				.clk(clk),
				.rstn(rstn),
				.a0(A0C80),
				.a1(A0C90),
				.a2(A0D80),
				.a3(A0D90),
				.p(P1640)
);

maxpool maxpool_47(
				.clk(clk),
				.rstn(rstn),
				.a0(A0CA0),
				.a1(A0CB0),
				.a2(A0DA0),
				.a3(A0DB0),
				.p(P1650)
);

maxpool maxpool_48(
				.clk(clk),
				.rstn(rstn),
				.a0(A0CC0),
				.a1(A0CD0),
				.a2(A0DC0),
				.a3(A0DD0),
				.p(P1660)
);

maxpool maxpool_49(
				.clk(clk),
				.rstn(rstn),
				.a0(A0001),
				.a1(A0011),
				.a2(A0101),
				.a3(A0111),
				.p(P1001)
);

maxpool maxpool_50(
				.clk(clk),
				.rstn(rstn),
				.a0(A0021),
				.a1(A0031),
				.a2(A0121),
				.a3(A0131),
				.p(P1011)
);

maxpool maxpool_51(
				.clk(clk),
				.rstn(rstn),
				.a0(A0041),
				.a1(A0051),
				.a2(A0141),
				.a3(A0151),
				.p(P1021)
);

maxpool maxpool_52(
				.clk(clk),
				.rstn(rstn),
				.a0(A0061),
				.a1(A0071),
				.a2(A0161),
				.a3(A0171),
				.p(P1031)
);

maxpool maxpool_53(
				.clk(clk),
				.rstn(rstn),
				.a0(A0081),
				.a1(A0091),
				.a2(A0181),
				.a3(A0191),
				.p(P1041)
);

maxpool maxpool_54(
				.clk(clk),
				.rstn(rstn),
				.a0(A00A1),
				.a1(A00B1),
				.a2(A01A1),
				.a3(A01B1),
				.p(P1051)
);

maxpool maxpool_55(
				.clk(clk),
				.rstn(rstn),
				.a0(A00C1),
				.a1(A00D1),
				.a2(A01C1),
				.a3(A01D1),
				.p(P1061)
);

maxpool maxpool_56(
				.clk(clk),
				.rstn(rstn),
				.a0(A0201),
				.a1(A0211),
				.a2(A0301),
				.a3(A0311),
				.p(P1101)
);

maxpool maxpool_57(
				.clk(clk),
				.rstn(rstn),
				.a0(A0221),
				.a1(A0231),
				.a2(A0321),
				.a3(A0331),
				.p(P1111)
);

maxpool maxpool_58(
				.clk(clk),
				.rstn(rstn),
				.a0(A0241),
				.a1(A0251),
				.a2(A0341),
				.a3(A0351),
				.p(P1121)
);

maxpool maxpool_59(
				.clk(clk),
				.rstn(rstn),
				.a0(A0261),
				.a1(A0271),
				.a2(A0361),
				.a3(A0371),
				.p(P1131)
);

maxpool maxpool_60(
				.clk(clk),
				.rstn(rstn),
				.a0(A0281),
				.a1(A0291),
				.a2(A0381),
				.a3(A0391),
				.p(P1141)
);

maxpool maxpool_61(
				.clk(clk),
				.rstn(rstn),
				.a0(A02A1),
				.a1(A02B1),
				.a2(A03A1),
				.a3(A03B1),
				.p(P1151)
);

maxpool maxpool_62(
				.clk(clk),
				.rstn(rstn),
				.a0(A02C1),
				.a1(A02D1),
				.a2(A03C1),
				.a3(A03D1),
				.p(P1161)
);

maxpool maxpool_63(
				.clk(clk),
				.rstn(rstn),
				.a0(A0401),
				.a1(A0411),
				.a2(A0501),
				.a3(A0511),
				.p(P1201)
);

maxpool maxpool_64(
				.clk(clk),
				.rstn(rstn),
				.a0(A0421),
				.a1(A0431),
				.a2(A0521),
				.a3(A0531),
				.p(P1211)
);

maxpool maxpool_65(
				.clk(clk),
				.rstn(rstn),
				.a0(A0441),
				.a1(A0451),
				.a2(A0541),
				.a3(A0551),
				.p(P1221)
);

maxpool maxpool_66(
				.clk(clk),
				.rstn(rstn),
				.a0(A0461),
				.a1(A0471),
				.a2(A0561),
				.a3(A0571),
				.p(P1231)
);

maxpool maxpool_67(
				.clk(clk),
				.rstn(rstn),
				.a0(A0481),
				.a1(A0491),
				.a2(A0581),
				.a3(A0591),
				.p(P1241)
);

maxpool maxpool_68(
				.clk(clk),
				.rstn(rstn),
				.a0(A04A1),
				.a1(A04B1),
				.a2(A05A1),
				.a3(A05B1),
				.p(P1251)
);

maxpool maxpool_69(
				.clk(clk),
				.rstn(rstn),
				.a0(A04C1),
				.a1(A04D1),
				.a2(A05C1),
				.a3(A05D1),
				.p(P1261)
);

maxpool maxpool_70(
				.clk(clk),
				.rstn(rstn),
				.a0(A0601),
				.a1(A0611),
				.a2(A0701),
				.a3(A0711),
				.p(P1301)
);

maxpool maxpool_71(
				.clk(clk),
				.rstn(rstn),
				.a0(A0621),
				.a1(A0631),
				.a2(A0721),
				.a3(A0731),
				.p(P1311)
);

maxpool maxpool_72(
				.clk(clk),
				.rstn(rstn),
				.a0(A0641),
				.a1(A0651),
				.a2(A0741),
				.a3(A0751),
				.p(P1321)
);

maxpool maxpool_73(
				.clk(clk),
				.rstn(rstn),
				.a0(A0661),
				.a1(A0671),
				.a2(A0761),
				.a3(A0771),
				.p(P1331)
);

maxpool maxpool_74(
				.clk(clk),
				.rstn(rstn),
				.a0(A0681),
				.a1(A0691),
				.a2(A0781),
				.a3(A0791),
				.p(P1341)
);

maxpool maxpool_75(
				.clk(clk),
				.rstn(rstn),
				.a0(A06A1),
				.a1(A06B1),
				.a2(A07A1),
				.a3(A07B1),
				.p(P1351)
);

maxpool maxpool_76(
				.clk(clk),
				.rstn(rstn),
				.a0(A06C1),
				.a1(A06D1),
				.a2(A07C1),
				.a3(A07D1),
				.p(P1361)
);

maxpool maxpool_77(
				.clk(clk),
				.rstn(rstn),
				.a0(A0801),
				.a1(A0811),
				.a2(A0901),
				.a3(A0911),
				.p(P1401)
);

maxpool maxpool_78(
				.clk(clk),
				.rstn(rstn),
				.a0(A0821),
				.a1(A0831),
				.a2(A0921),
				.a3(A0931),
				.p(P1411)
);

maxpool maxpool_79(
				.clk(clk),
				.rstn(rstn),
				.a0(A0841),
				.a1(A0851),
				.a2(A0941),
				.a3(A0951),
				.p(P1421)
);

maxpool maxpool_80(
				.clk(clk),
				.rstn(rstn),
				.a0(A0861),
				.a1(A0871),
				.a2(A0961),
				.a3(A0971),
				.p(P1431)
);

maxpool maxpool_81(
				.clk(clk),
				.rstn(rstn),
				.a0(A0881),
				.a1(A0891),
				.a2(A0981),
				.a3(A0991),
				.p(P1441)
);

maxpool maxpool_82(
				.clk(clk),
				.rstn(rstn),
				.a0(A08A1),
				.a1(A08B1),
				.a2(A09A1),
				.a3(A09B1),
				.p(P1451)
);

maxpool maxpool_83(
				.clk(clk),
				.rstn(rstn),
				.a0(A08C1),
				.a1(A08D1),
				.a2(A09C1),
				.a3(A09D1),
				.p(P1461)
);

maxpool maxpool_84(
				.clk(clk),
				.rstn(rstn),
				.a0(A0A01),
				.a1(A0A11),
				.a2(A0B01),
				.a3(A0B11),
				.p(P1501)
);

maxpool maxpool_85(
				.clk(clk),
				.rstn(rstn),
				.a0(A0A21),
				.a1(A0A31),
				.a2(A0B21),
				.a3(A0B31),
				.p(P1511)
);

maxpool maxpool_86(
				.clk(clk),
				.rstn(rstn),
				.a0(A0A41),
				.a1(A0A51),
				.a2(A0B41),
				.a3(A0B51),
				.p(P1521)
);

maxpool maxpool_87(
				.clk(clk),
				.rstn(rstn),
				.a0(A0A61),
				.a1(A0A71),
				.a2(A0B61),
				.a3(A0B71),
				.p(P1531)
);

maxpool maxpool_88(
				.clk(clk),
				.rstn(rstn),
				.a0(A0A81),
				.a1(A0A91),
				.a2(A0B81),
				.a3(A0B91),
				.p(P1541)
);

maxpool maxpool_89(
				.clk(clk),
				.rstn(rstn),
				.a0(A0AA1),
				.a1(A0AB1),
				.a2(A0BA1),
				.a3(A0BB1),
				.p(P1551)
);

maxpool maxpool_90(
				.clk(clk),
				.rstn(rstn),
				.a0(A0AC1),
				.a1(A0AD1),
				.a2(A0BC1),
				.a3(A0BD1),
				.p(P1561)
);

maxpool maxpool_91(
				.clk(clk),
				.rstn(rstn),
				.a0(A0C01),
				.a1(A0C11),
				.a2(A0D01),
				.a3(A0D11),
				.p(P1601)
);

maxpool maxpool_92(
				.clk(clk),
				.rstn(rstn),
				.a0(A0C21),
				.a1(A0C31),
				.a2(A0D21),
				.a3(A0D31),
				.p(P1611)
);

maxpool maxpool_93(
				.clk(clk),
				.rstn(rstn),
				.a0(A0C41),
				.a1(A0C51),
				.a2(A0D41),
				.a3(A0D51),
				.p(P1621)
);

maxpool maxpool_94(
				.clk(clk),
				.rstn(rstn),
				.a0(A0C61),
				.a1(A0C71),
				.a2(A0D61),
				.a3(A0D71),
				.p(P1631)
);

maxpool maxpool_95(
				.clk(clk),
				.rstn(rstn),
				.a0(A0C81),
				.a1(A0C91),
				.a2(A0D81),
				.a3(A0D91),
				.p(P1641)
);

maxpool maxpool_96(
				.clk(clk),
				.rstn(rstn),
				.a0(A0CA1),
				.a1(A0CB1),
				.a2(A0DA1),
				.a3(A0DB1),
				.p(P1651)
);

maxpool maxpool_97(
				.clk(clk),
				.rstn(rstn),
				.a0(A0CC1),
				.a1(A0CD1),
				.a2(A0DC1),
				.a3(A0DD1),
				.p(P1661)
);

maxpool maxpool_98(
				.clk(clk),
				.rstn(rstn),
				.a0(A0002),
				.a1(A0012),
				.a2(A0102),
				.a3(A0112),
				.p(P1002)
);

maxpool maxpool_99(
				.clk(clk),
				.rstn(rstn),
				.a0(A0022),
				.a1(A0032),
				.a2(A0122),
				.a3(A0132),
				.p(P1012)
);

maxpool maxpool_100(
				.clk(clk),
				.rstn(rstn),
				.a0(A0042),
				.a1(A0052),
				.a2(A0142),
				.a3(A0152),
				.p(P1022)
);

maxpool maxpool_101(
				.clk(clk),
				.rstn(rstn),
				.a0(A0062),
				.a1(A0072),
				.a2(A0162),
				.a3(A0172),
				.p(P1032)
);

maxpool maxpool_102(
				.clk(clk),
				.rstn(rstn),
				.a0(A0082),
				.a1(A0092),
				.a2(A0182),
				.a3(A0192),
				.p(P1042)
);

maxpool maxpool_103(
				.clk(clk),
				.rstn(rstn),
				.a0(A00A2),
				.a1(A00B2),
				.a2(A01A2),
				.a3(A01B2),
				.p(P1052)
);

maxpool maxpool_104(
				.clk(clk),
				.rstn(rstn),
				.a0(A00C2),
				.a1(A00D2),
				.a2(A01C2),
				.a3(A01D2),
				.p(P1062)
);

maxpool maxpool_105(
				.clk(clk),
				.rstn(rstn),
				.a0(A0202),
				.a1(A0212),
				.a2(A0302),
				.a3(A0312),
				.p(P1102)
);

maxpool maxpool_106(
				.clk(clk),
				.rstn(rstn),
				.a0(A0222),
				.a1(A0232),
				.a2(A0322),
				.a3(A0332),
				.p(P1112)
);

maxpool maxpool_107(
				.clk(clk),
				.rstn(rstn),
				.a0(A0242),
				.a1(A0252),
				.a2(A0342),
				.a3(A0352),
				.p(P1122)
);

maxpool maxpool_108(
				.clk(clk),
				.rstn(rstn),
				.a0(A0262),
				.a1(A0272),
				.a2(A0362),
				.a3(A0372),
				.p(P1132)
);

maxpool maxpool_109(
				.clk(clk),
				.rstn(rstn),
				.a0(A0282),
				.a1(A0292),
				.a2(A0382),
				.a3(A0392),
				.p(P1142)
);

maxpool maxpool_110(
				.clk(clk),
				.rstn(rstn),
				.a0(A02A2),
				.a1(A02B2),
				.a2(A03A2),
				.a3(A03B2),
				.p(P1152)
);

maxpool maxpool_111(
				.clk(clk),
				.rstn(rstn),
				.a0(A02C2),
				.a1(A02D2),
				.a2(A03C2),
				.a3(A03D2),
				.p(P1162)
);

maxpool maxpool_112(
				.clk(clk),
				.rstn(rstn),
				.a0(A0402),
				.a1(A0412),
				.a2(A0502),
				.a3(A0512),
				.p(P1202)
);

maxpool maxpool_113(
				.clk(clk),
				.rstn(rstn),
				.a0(A0422),
				.a1(A0432),
				.a2(A0522),
				.a3(A0532),
				.p(P1212)
);

maxpool maxpool_114(
				.clk(clk),
				.rstn(rstn),
				.a0(A0442),
				.a1(A0452),
				.a2(A0542),
				.a3(A0552),
				.p(P1222)
);

maxpool maxpool_115(
				.clk(clk),
				.rstn(rstn),
				.a0(A0462),
				.a1(A0472),
				.a2(A0562),
				.a3(A0572),
				.p(P1232)
);

maxpool maxpool_116(
				.clk(clk),
				.rstn(rstn),
				.a0(A0482),
				.a1(A0492),
				.a2(A0582),
				.a3(A0592),
				.p(P1242)
);

maxpool maxpool_117(
				.clk(clk),
				.rstn(rstn),
				.a0(A04A2),
				.a1(A04B2),
				.a2(A05A2),
				.a3(A05B2),
				.p(P1252)
);

maxpool maxpool_118(
				.clk(clk),
				.rstn(rstn),
				.a0(A04C2),
				.a1(A04D2),
				.a2(A05C2),
				.a3(A05D2),
				.p(P1262)
);

maxpool maxpool_119(
				.clk(clk),
				.rstn(rstn),
				.a0(A0602),
				.a1(A0612),
				.a2(A0702),
				.a3(A0712),
				.p(P1302)
);

maxpool maxpool_120(
				.clk(clk),
				.rstn(rstn),
				.a0(A0622),
				.a1(A0632),
				.a2(A0722),
				.a3(A0732),
				.p(P1312)
);

maxpool maxpool_121(
				.clk(clk),
				.rstn(rstn),
				.a0(A0642),
				.a1(A0652),
				.a2(A0742),
				.a3(A0752),
				.p(P1322)
);

maxpool maxpool_122(
				.clk(clk),
				.rstn(rstn),
				.a0(A0662),
				.a1(A0672),
				.a2(A0762),
				.a3(A0772),
				.p(P1332)
);

maxpool maxpool_123(
				.clk(clk),
				.rstn(rstn),
				.a0(A0682),
				.a1(A0692),
				.a2(A0782),
				.a3(A0792),
				.p(P1342)
);

maxpool maxpool_124(
				.clk(clk),
				.rstn(rstn),
				.a0(A06A2),
				.a1(A06B2),
				.a2(A07A2),
				.a3(A07B2),
				.p(P1352)
);

maxpool maxpool_125(
				.clk(clk),
				.rstn(rstn),
				.a0(A06C2),
				.a1(A06D2),
				.a2(A07C2),
				.a3(A07D2),
				.p(P1362)
);

maxpool maxpool_126(
				.clk(clk),
				.rstn(rstn),
				.a0(A0802),
				.a1(A0812),
				.a2(A0902),
				.a3(A0912),
				.p(P1402)
);

maxpool maxpool_127(
				.clk(clk),
				.rstn(rstn),
				.a0(A0822),
				.a1(A0832),
				.a2(A0922),
				.a3(A0932),
				.p(P1412)
);

maxpool maxpool_128(
				.clk(clk),
				.rstn(rstn),
				.a0(A0842),
				.a1(A0852),
				.a2(A0942),
				.a3(A0952),
				.p(P1422)
);

maxpool maxpool_129(
				.clk(clk),
				.rstn(rstn),
				.a0(A0862),
				.a1(A0872),
				.a2(A0962),
				.a3(A0972),
				.p(P1432)
);

maxpool maxpool_130(
				.clk(clk),
				.rstn(rstn),
				.a0(A0882),
				.a1(A0892),
				.a2(A0982),
				.a3(A0992),
				.p(P1442)
);

maxpool maxpool_131(
				.clk(clk),
				.rstn(rstn),
				.a0(A08A2),
				.a1(A08B2),
				.a2(A09A2),
				.a3(A09B2),
				.p(P1452)
);

maxpool maxpool_132(
				.clk(clk),
				.rstn(rstn),
				.a0(A08C2),
				.a1(A08D2),
				.a2(A09C2),
				.a3(A09D2),
				.p(P1462)
);

maxpool maxpool_133(
				.clk(clk),
				.rstn(rstn),
				.a0(A0A02),
				.a1(A0A12),
				.a2(A0B02),
				.a3(A0B12),
				.p(P1502)
);

maxpool maxpool_134(
				.clk(clk),
				.rstn(rstn),
				.a0(A0A22),
				.a1(A0A32),
				.a2(A0B22),
				.a3(A0B32),
				.p(P1512)
);

maxpool maxpool_135(
				.clk(clk),
				.rstn(rstn),
				.a0(A0A42),
				.a1(A0A52),
				.a2(A0B42),
				.a3(A0B52),
				.p(P1522)
);

maxpool maxpool_136(
				.clk(clk),
				.rstn(rstn),
				.a0(A0A62),
				.a1(A0A72),
				.a2(A0B62),
				.a3(A0B72),
				.p(P1532)
);

maxpool maxpool_137(
				.clk(clk),
				.rstn(rstn),
				.a0(A0A82),
				.a1(A0A92),
				.a2(A0B82),
				.a3(A0B92),
				.p(P1542)
);

maxpool maxpool_138(
				.clk(clk),
				.rstn(rstn),
				.a0(A0AA2),
				.a1(A0AB2),
				.a2(A0BA2),
				.a3(A0BB2),
				.p(P1552)
);

maxpool maxpool_139(
				.clk(clk),
				.rstn(rstn),
				.a0(A0AC2),
				.a1(A0AD2),
				.a2(A0BC2),
				.a3(A0BD2),
				.p(P1562)
);

maxpool maxpool_140(
				.clk(clk),
				.rstn(rstn),
				.a0(A0C02),
				.a1(A0C12),
				.a2(A0D02),
				.a3(A0D12),
				.p(P1602)
);

maxpool maxpool_141(
				.clk(clk),
				.rstn(rstn),
				.a0(A0C22),
				.a1(A0C32),
				.a2(A0D22),
				.a3(A0D32),
				.p(P1612)
);

maxpool maxpool_142(
				.clk(clk),
				.rstn(rstn),
				.a0(A0C42),
				.a1(A0C52),
				.a2(A0D42),
				.a3(A0D52),
				.p(P1622)
);

maxpool maxpool_143(
				.clk(clk),
				.rstn(rstn),
				.a0(A0C62),
				.a1(A0C72),
				.a2(A0D62),
				.a3(A0D72),
				.p(P1632)
);

maxpool maxpool_144(
				.clk(clk),
				.rstn(rstn),
				.a0(A0C82),
				.a1(A0C92),
				.a2(A0D82),
				.a3(A0D92),
				.p(P1642)
);

maxpool maxpool_145(
				.clk(clk),
				.rstn(rstn),
				.a0(A0CA2),
				.a1(A0CB2),
				.a2(A0DA2),
				.a3(A0DB2),
				.p(P1652)
);

maxpool maxpool_146(
				.clk(clk),
				.rstn(rstn),
				.a0(A0CC2),
				.a1(A0CD2),
				.a2(A0DC2),
				.a3(A0DD2),
				.p(P1662)
);

//layer1 done, begain next layer
wire P2000;
wire P2010;
wire P2020;
wire P2030;
wire P2040;
wire P2100;
wire P2110;
wire P2120;
wire P2130;
wire P2140;
wire P2200;
wire P2210;
wire P2220;
wire P2230;
wire P2240;
wire P2300;
wire P2310;
wire P2320;
wire P2330;
wire P2340;
wire P2400;
wire P2410;
wire P2420;
wire P2430;
wire P2440;
wire P2001;
wire P2011;
wire P2021;
wire P2031;
wire P2041;
wire P2101;
wire P2111;
wire P2121;
wire P2131;
wire P2141;
wire P2201;
wire P2211;
wire P2221;
wire P2231;
wire P2241;
wire P2301;
wire P2311;
wire P2321;
wire P2331;
wire P2341;
wire P2401;
wire P2411;
wire P2421;
wire P2431;
wire P2441;
wire P2002;
wire P2012;
wire P2022;
wire P2032;
wire P2042;
wire P2102;
wire P2112;
wire P2122;
wire P2132;
wire P2142;
wire P2202;
wire P2212;
wire P2222;
wire P2232;
wire P2242;
wire P2302;
wire P2312;
wire P2322;
wire P2332;
wire P2342;
wire P2402;
wire P2412;
wire P2422;
wire P2432;
wire P2442;
wire P2003;
wire P2013;
wire P2023;
wire P2033;
wire P2043;
wire P2103;
wire P2113;
wire P2123;
wire P2133;
wire P2143;
wire P2203;
wire P2213;
wire P2223;
wire P2233;
wire P2243;
wire P2303;
wire P2313;
wire P2323;
wire P2333;
wire P2343;
wire P2403;
wire P2413;
wire P2423;
wire P2433;
wire P2443;
wire P2004;
wire P2014;
wire P2024;
wire P2034;
wire P2044;
wire P2104;
wire P2114;
wire P2124;
wire P2134;
wire P2144;
wire P2204;
wire P2214;
wire P2224;
wire P2234;
wire P2244;
wire P2304;
wire P2314;
wire P2324;
wire P2334;
wire P2344;
wire P2404;
wire P2414;
wire P2424;
wire P2434;
wire P2444;
wire P2005;
wire P2015;
wire P2025;
wire P2035;
wire P2045;
wire P2105;
wire P2115;
wire P2125;
wire P2135;
wire P2145;
wire P2205;
wire P2215;
wire P2225;
wire P2235;
wire P2245;
wire P2305;
wire P2315;
wire P2325;
wire P2335;
wire P2345;
wire P2405;
wire P2415;
wire P2425;
wire P2435;
wire P2445;
wire P2006;
wire P2016;
wire P2026;
wire P2036;
wire P2046;
wire P2106;
wire P2116;
wire P2126;
wire P2136;
wire P2146;
wire P2206;
wire P2216;
wire P2226;
wire P2236;
wire P2246;
wire P2306;
wire P2316;
wire P2326;
wire P2336;
wire P2346;
wire P2406;
wire P2416;
wire P2426;
wire P2436;
wire P2446;
wire P2007;
wire P2017;
wire P2027;
wire P2037;
wire P2047;
wire P2107;
wire P2117;
wire P2127;
wire P2137;
wire P2147;
wire P2207;
wire P2217;
wire P2227;
wire P2237;
wire P2247;
wire P2307;
wire P2317;
wire P2327;
wire P2337;
wire P2347;
wire P2407;
wire P2417;
wire P2427;
wire P2437;
wire P2447;
wire P2008;
wire P2018;
wire P2028;
wire P2038;
wire P2048;
wire P2108;
wire P2118;
wire P2128;
wire P2138;
wire P2148;
wire P2208;
wire P2218;
wire P2228;
wire P2238;
wire P2248;
wire P2308;
wire P2318;
wire P2328;
wire P2338;
wire P2348;
wire P2408;
wire P2418;
wire P2428;
wire P2438;
wire P2448;
wire P2009;
wire P2019;
wire P2029;
wire P2039;
wire P2049;
wire P2109;
wire P2119;
wire P2129;
wire P2139;
wire P2149;
wire P2209;
wire P2219;
wire P2229;
wire P2239;
wire P2249;
wire P2309;
wire P2319;
wire P2329;
wire P2339;
wire P2349;
wire P2409;
wire P2419;
wire P2429;
wire P2439;
wire P2449;
wire P200A;
wire P201A;
wire P202A;
wire P203A;
wire P204A;
wire P210A;
wire P211A;
wire P212A;
wire P213A;
wire P214A;
wire P220A;
wire P221A;
wire P222A;
wire P223A;
wire P224A;
wire P230A;
wire P231A;
wire P232A;
wire P233A;
wire P234A;
wire P240A;
wire P241A;
wire P242A;
wire P243A;
wire P244A;
wire P200B;
wire P201B;
wire P202B;
wire P203B;
wire P204B;
wire P210B;
wire P211B;
wire P212B;
wire P213B;
wire P214B;
wire P220B;
wire P221B;
wire P222B;
wire P223B;
wire P224B;
wire P230B;
wire P231B;
wire P232B;
wire P233B;
wire P234B;
wire P240B;
wire P241B;
wire P242B;
wire P243B;
wire P244B;
wire P200C;
wire P201C;
wire P202C;
wire P203C;
wire P204C;
wire P210C;
wire P211C;
wire P212C;
wire P213C;
wire P214C;
wire P220C;
wire P221C;
wire P222C;
wire P223C;
wire P224C;
wire P230C;
wire P231C;
wire P232C;
wire P233C;
wire P234C;
wire P240C;
wire P241C;
wire P242C;
wire P243C;
wire P244C;
wire P200D;
wire P201D;
wire P202D;
wire P203D;
wire P204D;
wire P210D;
wire P211D;
wire P212D;
wire P213D;
wire P214D;
wire P220D;
wire P221D;
wire P222D;
wire P223D;
wire P224D;
wire P230D;
wire P231D;
wire P232D;
wire P233D;
wire P234D;
wire P240D;
wire P241D;
wire P242D;
wire P243D;
wire P244D;
wire P200E;
wire P201E;
wire P202E;
wire P203E;
wire P204E;
wire P210E;
wire P211E;
wire P212E;
wire P213E;
wire P214E;
wire P220E;
wire P221E;
wire P222E;
wire P223E;
wire P224E;
wire P230E;
wire P231E;
wire P232E;
wire P233E;
wire P234E;
wire P240E;
wire P241E;
wire P242E;
wire P243E;
wire P244E;
wire P200F;
wire P201F;
wire P202F;
wire P203F;
wire P204F;
wire P210F;
wire P211F;
wire P212F;
wire P213F;
wire P214F;
wire P220F;
wire P221F;
wire P222F;
wire P223F;
wire P224F;
wire P230F;
wire P231F;
wire P232F;
wire P233F;
wire P234F;
wire P240F;
wire P241F;
wire P242F;
wire P243F;
wire P244F;
wire W10000,W10010,W10020,W10100,W10110,W10120,W10200,W10210,W10220;
wire W10001,W10011,W10021,W10101,W10111,W10121,W10201,W10211,W10221;
wire W10002,W10012,W10022,W10102,W10112,W10122,W10202,W10212,W10222;
wire W11000,W11010,W11020,W11100,W11110,W11120,W11200,W11210,W11220;
wire W11001,W11011,W11021,W11101,W11111,W11121,W11201,W11211,W11221;
wire W11002,W11012,W11022,W11102,W11112,W11122,W11202,W11212,W11222;
wire W12000,W12010,W12020,W12100,W12110,W12120,W12200,W12210,W12220;
wire W12001,W12011,W12021,W12101,W12111,W12121,W12201,W12211,W12221;
wire W12002,W12012,W12022,W12102,W12112,W12122,W12202,W12212,W12222;
wire W13000,W13010,W13020,W13100,W13110,W13120,W13200,W13210,W13220;
wire W13001,W13011,W13021,W13101,W13111,W13121,W13201,W13211,W13221;
wire W13002,W13012,W13022,W13102,W13112,W13122,W13202,W13212,W13222;
wire W14000,W14010,W14020,W14100,W14110,W14120,W14200,W14210,W14220;
wire W14001,W14011,W14021,W14101,W14111,W14121,W14201,W14211,W14221;
wire W14002,W14012,W14022,W14102,W14112,W14122,W14202,W14212,W14222;
wire W15000,W15010,W15020,W15100,W15110,W15120,W15200,W15210,W15220;
wire W15001,W15011,W15021,W15101,W15111,W15121,W15201,W15211,W15221;
wire W15002,W15012,W15022,W15102,W15112,W15122,W15202,W15212,W15222;
wire W16000,W16010,W16020,W16100,W16110,W16120,W16200,W16210,W16220;
wire W16001,W16011,W16021,W16101,W16111,W16121,W16201,W16211,W16221;
wire W16002,W16012,W16022,W16102,W16112,W16122,W16202,W16212,W16222;
wire W17000,W17010,W17020,W17100,W17110,W17120,W17200,W17210,W17220;
wire W17001,W17011,W17021,W17101,W17111,W17121,W17201,W17211,W17221;
wire W17002,W17012,W17022,W17102,W17112,W17122,W17202,W17212,W17222;
wire W18000,W18010,W18020,W18100,W18110,W18120,W18200,W18210,W18220;
wire W18001,W18011,W18021,W18101,W18111,W18121,W18201,W18211,W18221;
wire W18002,W18012,W18022,W18102,W18112,W18122,W18202,W18212,W18222;
wire W19000,W19010,W19020,W19100,W19110,W19120,W19200,W19210,W19220;
wire W19001,W19011,W19021,W19101,W19111,W19121,W19201,W19211,W19221;
wire W19002,W19012,W19022,W19102,W19112,W19122,W19202,W19212,W19222;
wire W1A000,W1A010,W1A020,W1A100,W1A110,W1A120,W1A200,W1A210,W1A220;
wire W1A001,W1A011,W1A021,W1A101,W1A111,W1A121,W1A201,W1A211,W1A221;
wire W1A002,W1A012,W1A022,W1A102,W1A112,W1A122,W1A202,W1A212,W1A222;
wire W1B000,W1B010,W1B020,W1B100,W1B110,W1B120,W1B200,W1B210,W1B220;
wire W1B001,W1B011,W1B021,W1B101,W1B111,W1B121,W1B201,W1B211,W1B221;
wire W1B002,W1B012,W1B022,W1B102,W1B112,W1B122,W1B202,W1B212,W1B222;
wire W1C000,W1C010,W1C020,W1C100,W1C110,W1C120,W1C200,W1C210,W1C220;
wire W1C001,W1C011,W1C021,W1C101,W1C111,W1C121,W1C201,W1C211,W1C221;
wire W1C002,W1C012,W1C022,W1C102,W1C112,W1C122,W1C202,W1C212,W1C222;
wire W1D000,W1D010,W1D020,W1D100,W1D110,W1D120,W1D200,W1D210,W1D220;
wire W1D001,W1D011,W1D021,W1D101,W1D111,W1D121,W1D201,W1D211,W1D221;
wire W1D002,W1D012,W1D022,W1D102,W1D112,W1D122,W1D202,W1D212,W1D222;
wire W1E000,W1E010,W1E020,W1E100,W1E110,W1E120,W1E200,W1E210,W1E220;
wire W1E001,W1E011,W1E021,W1E101,W1E111,W1E121,W1E201,W1E211,W1E221;
wire W1E002,W1E012,W1E022,W1E102,W1E112,W1E122,W1E202,W1E212,W1E222;
wire W1F000,W1F010,W1F020,W1F100,W1F110,W1F120,W1F200,W1F210,W1F220;
wire W1F001,W1F011,W1F021,W1F101,W1F111,W1F121,W1F201,W1F211,W1F221;
wire W1F002,W1F012,W1F022,W1F102,W1F112,W1F122,W1F202,W1F212,W1F222;
wire signed [4:0] c10000,c11000,c12000;
wire signed [4:0] c10010,c11010,c12010;
wire signed [4:0] c10020,c11020,c12020;
wire signed [4:0] c10030,c11030,c12030;
wire signed [4:0] c10040,c11040,c12040;
wire signed [4:0] c10100,c11100,c12100;
wire signed [4:0] c10110,c11110,c12110;
wire signed [4:0] c10120,c11120,c12120;
wire signed [4:0] c10130,c11130,c12130;
wire signed [4:0] c10140,c11140,c12140;
wire signed [4:0] c10200,c11200,c12200;
wire signed [4:0] c10210,c11210,c12210;
wire signed [4:0] c10220,c11220,c12220;
wire signed [4:0] c10230,c11230,c12230;
wire signed [4:0] c10240,c11240,c12240;
wire signed [4:0] c10300,c11300,c12300;
wire signed [4:0] c10310,c11310,c12310;
wire signed [4:0] c10320,c11320,c12320;
wire signed [4:0] c10330,c11330,c12330;
wire signed [4:0] c10340,c11340,c12340;
wire signed [4:0] c10400,c11400,c12400;
wire signed [4:0] c10410,c11410,c12410;
wire signed [4:0] c10420,c11420,c12420;
wire signed [4:0] c10430,c11430,c12430;
wire signed [4:0] c10440,c11440,c12440;
wire signed [4:0] c10001,c11001,c12001;
wire signed [4:0] c10011,c11011,c12011;
wire signed [4:0] c10021,c11021,c12021;
wire signed [4:0] c10031,c11031,c12031;
wire signed [4:0] c10041,c11041,c12041;
wire signed [4:0] c10101,c11101,c12101;
wire signed [4:0] c10111,c11111,c12111;
wire signed [4:0] c10121,c11121,c12121;
wire signed [4:0] c10131,c11131,c12131;
wire signed [4:0] c10141,c11141,c12141;
wire signed [4:0] c10201,c11201,c12201;
wire signed [4:0] c10211,c11211,c12211;
wire signed [4:0] c10221,c11221,c12221;
wire signed [4:0] c10231,c11231,c12231;
wire signed [4:0] c10241,c11241,c12241;
wire signed [4:0] c10301,c11301,c12301;
wire signed [4:0] c10311,c11311,c12311;
wire signed [4:0] c10321,c11321,c12321;
wire signed [4:0] c10331,c11331,c12331;
wire signed [4:0] c10341,c11341,c12341;
wire signed [4:0] c10401,c11401,c12401;
wire signed [4:0] c10411,c11411,c12411;
wire signed [4:0] c10421,c11421,c12421;
wire signed [4:0] c10431,c11431,c12431;
wire signed [4:0] c10441,c11441,c12441;
wire signed [4:0] c10002,c11002,c12002;
wire signed [4:0] c10012,c11012,c12012;
wire signed [4:0] c10022,c11022,c12022;
wire signed [4:0] c10032,c11032,c12032;
wire signed [4:0] c10042,c11042,c12042;
wire signed [4:0] c10102,c11102,c12102;
wire signed [4:0] c10112,c11112,c12112;
wire signed [4:0] c10122,c11122,c12122;
wire signed [4:0] c10132,c11132,c12132;
wire signed [4:0] c10142,c11142,c12142;
wire signed [4:0] c10202,c11202,c12202;
wire signed [4:0] c10212,c11212,c12212;
wire signed [4:0] c10222,c11222,c12222;
wire signed [4:0] c10232,c11232,c12232;
wire signed [4:0] c10242,c11242,c12242;
wire signed [4:0] c10302,c11302,c12302;
wire signed [4:0] c10312,c11312,c12312;
wire signed [4:0] c10322,c11322,c12322;
wire signed [4:0] c10332,c11332,c12332;
wire signed [4:0] c10342,c11342,c12342;
wire signed [4:0] c10402,c11402,c12402;
wire signed [4:0] c10412,c11412,c12412;
wire signed [4:0] c10422,c11422,c12422;
wire signed [4:0] c10432,c11432,c12432;
wire signed [4:0] c10442,c11442,c12442;
wire signed [4:0] c10003,c11003,c12003;
wire signed [4:0] c10013,c11013,c12013;
wire signed [4:0] c10023,c11023,c12023;
wire signed [4:0] c10033,c11033,c12033;
wire signed [4:0] c10043,c11043,c12043;
wire signed [4:0] c10103,c11103,c12103;
wire signed [4:0] c10113,c11113,c12113;
wire signed [4:0] c10123,c11123,c12123;
wire signed [4:0] c10133,c11133,c12133;
wire signed [4:0] c10143,c11143,c12143;
wire signed [4:0] c10203,c11203,c12203;
wire signed [4:0] c10213,c11213,c12213;
wire signed [4:0] c10223,c11223,c12223;
wire signed [4:0] c10233,c11233,c12233;
wire signed [4:0] c10243,c11243,c12243;
wire signed [4:0] c10303,c11303,c12303;
wire signed [4:0] c10313,c11313,c12313;
wire signed [4:0] c10323,c11323,c12323;
wire signed [4:0] c10333,c11333,c12333;
wire signed [4:0] c10343,c11343,c12343;
wire signed [4:0] c10403,c11403,c12403;
wire signed [4:0] c10413,c11413,c12413;
wire signed [4:0] c10423,c11423,c12423;
wire signed [4:0] c10433,c11433,c12433;
wire signed [4:0] c10443,c11443,c12443;
wire signed [4:0] c10004,c11004,c12004;
wire signed [4:0] c10014,c11014,c12014;
wire signed [4:0] c10024,c11024,c12024;
wire signed [4:0] c10034,c11034,c12034;
wire signed [4:0] c10044,c11044,c12044;
wire signed [4:0] c10104,c11104,c12104;
wire signed [4:0] c10114,c11114,c12114;
wire signed [4:0] c10124,c11124,c12124;
wire signed [4:0] c10134,c11134,c12134;
wire signed [4:0] c10144,c11144,c12144;
wire signed [4:0] c10204,c11204,c12204;
wire signed [4:0] c10214,c11214,c12214;
wire signed [4:0] c10224,c11224,c12224;
wire signed [4:0] c10234,c11234,c12234;
wire signed [4:0] c10244,c11244,c12244;
wire signed [4:0] c10304,c11304,c12304;
wire signed [4:0] c10314,c11314,c12314;
wire signed [4:0] c10324,c11324,c12324;
wire signed [4:0] c10334,c11334,c12334;
wire signed [4:0] c10344,c11344,c12344;
wire signed [4:0] c10404,c11404,c12404;
wire signed [4:0] c10414,c11414,c12414;
wire signed [4:0] c10424,c11424,c12424;
wire signed [4:0] c10434,c11434,c12434;
wire signed [4:0] c10444,c11444,c12444;
wire signed [4:0] c10005,c11005,c12005;
wire signed [4:0] c10015,c11015,c12015;
wire signed [4:0] c10025,c11025,c12025;
wire signed [4:0] c10035,c11035,c12035;
wire signed [4:0] c10045,c11045,c12045;
wire signed [4:0] c10105,c11105,c12105;
wire signed [4:0] c10115,c11115,c12115;
wire signed [4:0] c10125,c11125,c12125;
wire signed [4:0] c10135,c11135,c12135;
wire signed [4:0] c10145,c11145,c12145;
wire signed [4:0] c10205,c11205,c12205;
wire signed [4:0] c10215,c11215,c12215;
wire signed [4:0] c10225,c11225,c12225;
wire signed [4:0] c10235,c11235,c12235;
wire signed [4:0] c10245,c11245,c12245;
wire signed [4:0] c10305,c11305,c12305;
wire signed [4:0] c10315,c11315,c12315;
wire signed [4:0] c10325,c11325,c12325;
wire signed [4:0] c10335,c11335,c12335;
wire signed [4:0] c10345,c11345,c12345;
wire signed [4:0] c10405,c11405,c12405;
wire signed [4:0] c10415,c11415,c12415;
wire signed [4:0] c10425,c11425,c12425;
wire signed [4:0] c10435,c11435,c12435;
wire signed [4:0] c10445,c11445,c12445;
wire signed [4:0] c10006,c11006,c12006;
wire signed [4:0] c10016,c11016,c12016;
wire signed [4:0] c10026,c11026,c12026;
wire signed [4:0] c10036,c11036,c12036;
wire signed [4:0] c10046,c11046,c12046;
wire signed [4:0] c10106,c11106,c12106;
wire signed [4:0] c10116,c11116,c12116;
wire signed [4:0] c10126,c11126,c12126;
wire signed [4:0] c10136,c11136,c12136;
wire signed [4:0] c10146,c11146,c12146;
wire signed [4:0] c10206,c11206,c12206;
wire signed [4:0] c10216,c11216,c12216;
wire signed [4:0] c10226,c11226,c12226;
wire signed [4:0] c10236,c11236,c12236;
wire signed [4:0] c10246,c11246,c12246;
wire signed [4:0] c10306,c11306,c12306;
wire signed [4:0] c10316,c11316,c12316;
wire signed [4:0] c10326,c11326,c12326;
wire signed [4:0] c10336,c11336,c12336;
wire signed [4:0] c10346,c11346,c12346;
wire signed [4:0] c10406,c11406,c12406;
wire signed [4:0] c10416,c11416,c12416;
wire signed [4:0] c10426,c11426,c12426;
wire signed [4:0] c10436,c11436,c12436;
wire signed [4:0] c10446,c11446,c12446;
wire signed [4:0] c10007,c11007,c12007;
wire signed [4:0] c10017,c11017,c12017;
wire signed [4:0] c10027,c11027,c12027;
wire signed [4:0] c10037,c11037,c12037;
wire signed [4:0] c10047,c11047,c12047;
wire signed [4:0] c10107,c11107,c12107;
wire signed [4:0] c10117,c11117,c12117;
wire signed [4:0] c10127,c11127,c12127;
wire signed [4:0] c10137,c11137,c12137;
wire signed [4:0] c10147,c11147,c12147;
wire signed [4:0] c10207,c11207,c12207;
wire signed [4:0] c10217,c11217,c12217;
wire signed [4:0] c10227,c11227,c12227;
wire signed [4:0] c10237,c11237,c12237;
wire signed [4:0] c10247,c11247,c12247;
wire signed [4:0] c10307,c11307,c12307;
wire signed [4:0] c10317,c11317,c12317;
wire signed [4:0] c10327,c11327,c12327;
wire signed [4:0] c10337,c11337,c12337;
wire signed [4:0] c10347,c11347,c12347;
wire signed [4:0] c10407,c11407,c12407;
wire signed [4:0] c10417,c11417,c12417;
wire signed [4:0] c10427,c11427,c12427;
wire signed [4:0] c10437,c11437,c12437;
wire signed [4:0] c10447,c11447,c12447;
wire signed [4:0] c10008,c11008,c12008;
wire signed [4:0] c10018,c11018,c12018;
wire signed [4:0] c10028,c11028,c12028;
wire signed [4:0] c10038,c11038,c12038;
wire signed [4:0] c10048,c11048,c12048;
wire signed [4:0] c10108,c11108,c12108;
wire signed [4:0] c10118,c11118,c12118;
wire signed [4:0] c10128,c11128,c12128;
wire signed [4:0] c10138,c11138,c12138;
wire signed [4:0] c10148,c11148,c12148;
wire signed [4:0] c10208,c11208,c12208;
wire signed [4:0] c10218,c11218,c12218;
wire signed [4:0] c10228,c11228,c12228;
wire signed [4:0] c10238,c11238,c12238;
wire signed [4:0] c10248,c11248,c12248;
wire signed [4:0] c10308,c11308,c12308;
wire signed [4:0] c10318,c11318,c12318;
wire signed [4:0] c10328,c11328,c12328;
wire signed [4:0] c10338,c11338,c12338;
wire signed [4:0] c10348,c11348,c12348;
wire signed [4:0] c10408,c11408,c12408;
wire signed [4:0] c10418,c11418,c12418;
wire signed [4:0] c10428,c11428,c12428;
wire signed [4:0] c10438,c11438,c12438;
wire signed [4:0] c10448,c11448,c12448;
wire signed [4:0] c10009,c11009,c12009;
wire signed [4:0] c10019,c11019,c12019;
wire signed [4:0] c10029,c11029,c12029;
wire signed [4:0] c10039,c11039,c12039;
wire signed [4:0] c10049,c11049,c12049;
wire signed [4:0] c10109,c11109,c12109;
wire signed [4:0] c10119,c11119,c12119;
wire signed [4:0] c10129,c11129,c12129;
wire signed [4:0] c10139,c11139,c12139;
wire signed [4:0] c10149,c11149,c12149;
wire signed [4:0] c10209,c11209,c12209;
wire signed [4:0] c10219,c11219,c12219;
wire signed [4:0] c10229,c11229,c12229;
wire signed [4:0] c10239,c11239,c12239;
wire signed [4:0] c10249,c11249,c12249;
wire signed [4:0] c10309,c11309,c12309;
wire signed [4:0] c10319,c11319,c12319;
wire signed [4:0] c10329,c11329,c12329;
wire signed [4:0] c10339,c11339,c12339;
wire signed [4:0] c10349,c11349,c12349;
wire signed [4:0] c10409,c11409,c12409;
wire signed [4:0] c10419,c11419,c12419;
wire signed [4:0] c10429,c11429,c12429;
wire signed [4:0] c10439,c11439,c12439;
wire signed [4:0] c10449,c11449,c12449;
wire signed [4:0] c1000A,c1100A,c1200A;
wire signed [4:0] c1001A,c1101A,c1201A;
wire signed [4:0] c1002A,c1102A,c1202A;
wire signed [4:0] c1003A,c1103A,c1203A;
wire signed [4:0] c1004A,c1104A,c1204A;
wire signed [4:0] c1010A,c1110A,c1210A;
wire signed [4:0] c1011A,c1111A,c1211A;
wire signed [4:0] c1012A,c1112A,c1212A;
wire signed [4:0] c1013A,c1113A,c1213A;
wire signed [4:0] c1014A,c1114A,c1214A;
wire signed [4:0] c1020A,c1120A,c1220A;
wire signed [4:0] c1021A,c1121A,c1221A;
wire signed [4:0] c1022A,c1122A,c1222A;
wire signed [4:0] c1023A,c1123A,c1223A;
wire signed [4:0] c1024A,c1124A,c1224A;
wire signed [4:0] c1030A,c1130A,c1230A;
wire signed [4:0] c1031A,c1131A,c1231A;
wire signed [4:0] c1032A,c1132A,c1232A;
wire signed [4:0] c1033A,c1133A,c1233A;
wire signed [4:0] c1034A,c1134A,c1234A;
wire signed [4:0] c1040A,c1140A,c1240A;
wire signed [4:0] c1041A,c1141A,c1241A;
wire signed [4:0] c1042A,c1142A,c1242A;
wire signed [4:0] c1043A,c1143A,c1243A;
wire signed [4:0] c1044A,c1144A,c1244A;
wire signed [4:0] c1000B,c1100B,c1200B;
wire signed [4:0] c1001B,c1101B,c1201B;
wire signed [4:0] c1002B,c1102B,c1202B;
wire signed [4:0] c1003B,c1103B,c1203B;
wire signed [4:0] c1004B,c1104B,c1204B;
wire signed [4:0] c1010B,c1110B,c1210B;
wire signed [4:0] c1011B,c1111B,c1211B;
wire signed [4:0] c1012B,c1112B,c1212B;
wire signed [4:0] c1013B,c1113B,c1213B;
wire signed [4:0] c1014B,c1114B,c1214B;
wire signed [4:0] c1020B,c1120B,c1220B;
wire signed [4:0] c1021B,c1121B,c1221B;
wire signed [4:0] c1022B,c1122B,c1222B;
wire signed [4:0] c1023B,c1123B,c1223B;
wire signed [4:0] c1024B,c1124B,c1224B;
wire signed [4:0] c1030B,c1130B,c1230B;
wire signed [4:0] c1031B,c1131B,c1231B;
wire signed [4:0] c1032B,c1132B,c1232B;
wire signed [4:0] c1033B,c1133B,c1233B;
wire signed [4:0] c1034B,c1134B,c1234B;
wire signed [4:0] c1040B,c1140B,c1240B;
wire signed [4:0] c1041B,c1141B,c1241B;
wire signed [4:0] c1042B,c1142B,c1242B;
wire signed [4:0] c1043B,c1143B,c1243B;
wire signed [4:0] c1044B,c1144B,c1244B;
wire signed [4:0] c1000C,c1100C,c1200C;
wire signed [4:0] c1001C,c1101C,c1201C;
wire signed [4:0] c1002C,c1102C,c1202C;
wire signed [4:0] c1003C,c1103C,c1203C;
wire signed [4:0] c1004C,c1104C,c1204C;
wire signed [4:0] c1010C,c1110C,c1210C;
wire signed [4:0] c1011C,c1111C,c1211C;
wire signed [4:0] c1012C,c1112C,c1212C;
wire signed [4:0] c1013C,c1113C,c1213C;
wire signed [4:0] c1014C,c1114C,c1214C;
wire signed [4:0] c1020C,c1120C,c1220C;
wire signed [4:0] c1021C,c1121C,c1221C;
wire signed [4:0] c1022C,c1122C,c1222C;
wire signed [4:0] c1023C,c1123C,c1223C;
wire signed [4:0] c1024C,c1124C,c1224C;
wire signed [4:0] c1030C,c1130C,c1230C;
wire signed [4:0] c1031C,c1131C,c1231C;
wire signed [4:0] c1032C,c1132C,c1232C;
wire signed [4:0] c1033C,c1133C,c1233C;
wire signed [4:0] c1034C,c1134C,c1234C;
wire signed [4:0] c1040C,c1140C,c1240C;
wire signed [4:0] c1041C,c1141C,c1241C;
wire signed [4:0] c1042C,c1142C,c1242C;
wire signed [4:0] c1043C,c1143C,c1243C;
wire signed [4:0] c1044C,c1144C,c1244C;
wire signed [4:0] c1000D,c1100D,c1200D;
wire signed [4:0] c1001D,c1101D,c1201D;
wire signed [4:0] c1002D,c1102D,c1202D;
wire signed [4:0] c1003D,c1103D,c1203D;
wire signed [4:0] c1004D,c1104D,c1204D;
wire signed [4:0] c1010D,c1110D,c1210D;
wire signed [4:0] c1011D,c1111D,c1211D;
wire signed [4:0] c1012D,c1112D,c1212D;
wire signed [4:0] c1013D,c1113D,c1213D;
wire signed [4:0] c1014D,c1114D,c1214D;
wire signed [4:0] c1020D,c1120D,c1220D;
wire signed [4:0] c1021D,c1121D,c1221D;
wire signed [4:0] c1022D,c1122D,c1222D;
wire signed [4:0] c1023D,c1123D,c1223D;
wire signed [4:0] c1024D,c1124D,c1224D;
wire signed [4:0] c1030D,c1130D,c1230D;
wire signed [4:0] c1031D,c1131D,c1231D;
wire signed [4:0] c1032D,c1132D,c1232D;
wire signed [4:0] c1033D,c1133D,c1233D;
wire signed [4:0] c1034D,c1134D,c1234D;
wire signed [4:0] c1040D,c1140D,c1240D;
wire signed [4:0] c1041D,c1141D,c1241D;
wire signed [4:0] c1042D,c1142D,c1242D;
wire signed [4:0] c1043D,c1143D,c1243D;
wire signed [4:0] c1044D,c1144D,c1244D;
wire signed [4:0] c1000E,c1100E,c1200E;
wire signed [4:0] c1001E,c1101E,c1201E;
wire signed [4:0] c1002E,c1102E,c1202E;
wire signed [4:0] c1003E,c1103E,c1203E;
wire signed [4:0] c1004E,c1104E,c1204E;
wire signed [4:0] c1010E,c1110E,c1210E;
wire signed [4:0] c1011E,c1111E,c1211E;
wire signed [4:0] c1012E,c1112E,c1212E;
wire signed [4:0] c1013E,c1113E,c1213E;
wire signed [4:0] c1014E,c1114E,c1214E;
wire signed [4:0] c1020E,c1120E,c1220E;
wire signed [4:0] c1021E,c1121E,c1221E;
wire signed [4:0] c1022E,c1122E,c1222E;
wire signed [4:0] c1023E,c1123E,c1223E;
wire signed [4:0] c1024E,c1124E,c1224E;
wire signed [4:0] c1030E,c1130E,c1230E;
wire signed [4:0] c1031E,c1131E,c1231E;
wire signed [4:0] c1032E,c1132E,c1232E;
wire signed [4:0] c1033E,c1133E,c1233E;
wire signed [4:0] c1034E,c1134E,c1234E;
wire signed [4:0] c1040E,c1140E,c1240E;
wire signed [4:0] c1041E,c1141E,c1241E;
wire signed [4:0] c1042E,c1142E,c1242E;
wire signed [4:0] c1043E,c1143E,c1243E;
wire signed [4:0] c1044E,c1144E,c1244E;
wire signed [4:0] c1000F,c1100F,c1200F;
wire signed [4:0] c1001F,c1101F,c1201F;
wire signed [4:0] c1002F,c1102F,c1202F;
wire signed [4:0] c1003F,c1103F,c1203F;
wire signed [4:0] c1004F,c1104F,c1204F;
wire signed [4:0] c1010F,c1110F,c1210F;
wire signed [4:0] c1011F,c1111F,c1211F;
wire signed [4:0] c1012F,c1112F,c1212F;
wire signed [4:0] c1013F,c1113F,c1213F;
wire signed [4:0] c1014F,c1114F,c1214F;
wire signed [4:0] c1020F,c1120F,c1220F;
wire signed [4:0] c1021F,c1121F,c1221F;
wire signed [4:0] c1022F,c1122F,c1222F;
wire signed [4:0] c1023F,c1123F,c1223F;
wire signed [4:0] c1024F,c1124F,c1224F;
wire signed [4:0] c1030F,c1130F,c1230F;
wire signed [4:0] c1031F,c1131F,c1231F;
wire signed [4:0] c1032F,c1132F,c1232F;
wire signed [4:0] c1033F,c1133F,c1233F;
wire signed [4:0] c1034F,c1134F,c1234F;
wire signed [4:0] c1040F,c1140F,c1240F;
wire signed [4:0] c1041F,c1141F,c1241F;
wire signed [4:0] c1042F,c1142F,c1242F;
wire signed [4:0] c1043F,c1143F,c1243F;
wire signed [4:0] c1044F,c1144F,c1244F;
wire signed [6:0] C1000;
wire A1000;
wire signed [6:0] C1010;
wire A1010;
wire signed [6:0] C1020;
wire A1020;
wire signed [6:0] C1030;
wire A1030;
wire signed [6:0] C1040;
wire A1040;
wire signed [6:0] C1100;
wire A1100;
wire signed [6:0] C1110;
wire A1110;
wire signed [6:0] C1120;
wire A1120;
wire signed [6:0] C1130;
wire A1130;
wire signed [6:0] C1140;
wire A1140;
wire signed [6:0] C1200;
wire A1200;
wire signed [6:0] C1210;
wire A1210;
wire signed [6:0] C1220;
wire A1220;
wire signed [6:0] C1230;
wire A1230;
wire signed [6:0] C1240;
wire A1240;
wire signed [6:0] C1300;
wire A1300;
wire signed [6:0] C1310;
wire A1310;
wire signed [6:0] C1320;
wire A1320;
wire signed [6:0] C1330;
wire A1330;
wire signed [6:0] C1340;
wire A1340;
wire signed [6:0] C1400;
wire A1400;
wire signed [6:0] C1410;
wire A1410;
wire signed [6:0] C1420;
wire A1420;
wire signed [6:0] C1430;
wire A1430;
wire signed [6:0] C1440;
wire A1440;
wire signed [6:0] C1001;
wire A1001;
wire signed [6:0] C1011;
wire A1011;
wire signed [6:0] C1021;
wire A1021;
wire signed [6:0] C1031;
wire A1031;
wire signed [6:0] C1041;
wire A1041;
wire signed [6:0] C1101;
wire A1101;
wire signed [6:0] C1111;
wire A1111;
wire signed [6:0] C1121;
wire A1121;
wire signed [6:0] C1131;
wire A1131;
wire signed [6:0] C1141;
wire A1141;
wire signed [6:0] C1201;
wire A1201;
wire signed [6:0] C1211;
wire A1211;
wire signed [6:0] C1221;
wire A1221;
wire signed [6:0] C1231;
wire A1231;
wire signed [6:0] C1241;
wire A1241;
wire signed [6:0] C1301;
wire A1301;
wire signed [6:0] C1311;
wire A1311;
wire signed [6:0] C1321;
wire A1321;
wire signed [6:0] C1331;
wire A1331;
wire signed [6:0] C1341;
wire A1341;
wire signed [6:0] C1401;
wire A1401;
wire signed [6:0] C1411;
wire A1411;
wire signed [6:0] C1421;
wire A1421;
wire signed [6:0] C1431;
wire A1431;
wire signed [6:0] C1441;
wire A1441;
wire signed [6:0] C1002;
wire A1002;
wire signed [6:0] C1012;
wire A1012;
wire signed [6:0] C1022;
wire A1022;
wire signed [6:0] C1032;
wire A1032;
wire signed [6:0] C1042;
wire A1042;
wire signed [6:0] C1102;
wire A1102;
wire signed [6:0] C1112;
wire A1112;
wire signed [6:0] C1122;
wire A1122;
wire signed [6:0] C1132;
wire A1132;
wire signed [6:0] C1142;
wire A1142;
wire signed [6:0] C1202;
wire A1202;
wire signed [6:0] C1212;
wire A1212;
wire signed [6:0] C1222;
wire A1222;
wire signed [6:0] C1232;
wire A1232;
wire signed [6:0] C1242;
wire A1242;
wire signed [6:0] C1302;
wire A1302;
wire signed [6:0] C1312;
wire A1312;
wire signed [6:0] C1322;
wire A1322;
wire signed [6:0] C1332;
wire A1332;
wire signed [6:0] C1342;
wire A1342;
wire signed [6:0] C1402;
wire A1402;
wire signed [6:0] C1412;
wire A1412;
wire signed [6:0] C1422;
wire A1422;
wire signed [6:0] C1432;
wire A1432;
wire signed [6:0] C1442;
wire A1442;
wire signed [6:0] C1003;
wire A1003;
wire signed [6:0] C1013;
wire A1013;
wire signed [6:0] C1023;
wire A1023;
wire signed [6:0] C1033;
wire A1033;
wire signed [6:0] C1043;
wire A1043;
wire signed [6:0] C1103;
wire A1103;
wire signed [6:0] C1113;
wire A1113;
wire signed [6:0] C1123;
wire A1123;
wire signed [6:0] C1133;
wire A1133;
wire signed [6:0] C1143;
wire A1143;
wire signed [6:0] C1203;
wire A1203;
wire signed [6:0] C1213;
wire A1213;
wire signed [6:0] C1223;
wire A1223;
wire signed [6:0] C1233;
wire A1233;
wire signed [6:0] C1243;
wire A1243;
wire signed [6:0] C1303;
wire A1303;
wire signed [6:0] C1313;
wire A1313;
wire signed [6:0] C1323;
wire A1323;
wire signed [6:0] C1333;
wire A1333;
wire signed [6:0] C1343;
wire A1343;
wire signed [6:0] C1403;
wire A1403;
wire signed [6:0] C1413;
wire A1413;
wire signed [6:0] C1423;
wire A1423;
wire signed [6:0] C1433;
wire A1433;
wire signed [6:0] C1443;
wire A1443;
wire signed [6:0] C1004;
wire A1004;
wire signed [6:0] C1014;
wire A1014;
wire signed [6:0] C1024;
wire A1024;
wire signed [6:0] C1034;
wire A1034;
wire signed [6:0] C1044;
wire A1044;
wire signed [6:0] C1104;
wire A1104;
wire signed [6:0] C1114;
wire A1114;
wire signed [6:0] C1124;
wire A1124;
wire signed [6:0] C1134;
wire A1134;
wire signed [6:0] C1144;
wire A1144;
wire signed [6:0] C1204;
wire A1204;
wire signed [6:0] C1214;
wire A1214;
wire signed [6:0] C1224;
wire A1224;
wire signed [6:0] C1234;
wire A1234;
wire signed [6:0] C1244;
wire A1244;
wire signed [6:0] C1304;
wire A1304;
wire signed [6:0] C1314;
wire A1314;
wire signed [6:0] C1324;
wire A1324;
wire signed [6:0] C1334;
wire A1334;
wire signed [6:0] C1344;
wire A1344;
wire signed [6:0] C1404;
wire A1404;
wire signed [6:0] C1414;
wire A1414;
wire signed [6:0] C1424;
wire A1424;
wire signed [6:0] C1434;
wire A1434;
wire signed [6:0] C1444;
wire A1444;
wire signed [6:0] C1005;
wire A1005;
wire signed [6:0] C1015;
wire A1015;
wire signed [6:0] C1025;
wire A1025;
wire signed [6:0] C1035;
wire A1035;
wire signed [6:0] C1045;
wire A1045;
wire signed [6:0] C1105;
wire A1105;
wire signed [6:0] C1115;
wire A1115;
wire signed [6:0] C1125;
wire A1125;
wire signed [6:0] C1135;
wire A1135;
wire signed [6:0] C1145;
wire A1145;
wire signed [6:0] C1205;
wire A1205;
wire signed [6:0] C1215;
wire A1215;
wire signed [6:0] C1225;
wire A1225;
wire signed [6:0] C1235;
wire A1235;
wire signed [6:0] C1245;
wire A1245;
wire signed [6:0] C1305;
wire A1305;
wire signed [6:0] C1315;
wire A1315;
wire signed [6:0] C1325;
wire A1325;
wire signed [6:0] C1335;
wire A1335;
wire signed [6:0] C1345;
wire A1345;
wire signed [6:0] C1405;
wire A1405;
wire signed [6:0] C1415;
wire A1415;
wire signed [6:0] C1425;
wire A1425;
wire signed [6:0] C1435;
wire A1435;
wire signed [6:0] C1445;
wire A1445;
wire signed [6:0] C1006;
wire A1006;
wire signed [6:0] C1016;
wire A1016;
wire signed [6:0] C1026;
wire A1026;
wire signed [6:0] C1036;
wire A1036;
wire signed [6:0] C1046;
wire A1046;
wire signed [6:0] C1106;
wire A1106;
wire signed [6:0] C1116;
wire A1116;
wire signed [6:0] C1126;
wire A1126;
wire signed [6:0] C1136;
wire A1136;
wire signed [6:0] C1146;
wire A1146;
wire signed [6:0] C1206;
wire A1206;
wire signed [6:0] C1216;
wire A1216;
wire signed [6:0] C1226;
wire A1226;
wire signed [6:0] C1236;
wire A1236;
wire signed [6:0] C1246;
wire A1246;
wire signed [6:0] C1306;
wire A1306;
wire signed [6:0] C1316;
wire A1316;
wire signed [6:0] C1326;
wire A1326;
wire signed [6:0] C1336;
wire A1336;
wire signed [6:0] C1346;
wire A1346;
wire signed [6:0] C1406;
wire A1406;
wire signed [6:0] C1416;
wire A1416;
wire signed [6:0] C1426;
wire A1426;
wire signed [6:0] C1436;
wire A1436;
wire signed [6:0] C1446;
wire A1446;
wire signed [6:0] C1007;
wire A1007;
wire signed [6:0] C1017;
wire A1017;
wire signed [6:0] C1027;
wire A1027;
wire signed [6:0] C1037;
wire A1037;
wire signed [6:0] C1047;
wire A1047;
wire signed [6:0] C1107;
wire A1107;
wire signed [6:0] C1117;
wire A1117;
wire signed [6:0] C1127;
wire A1127;
wire signed [6:0] C1137;
wire A1137;
wire signed [6:0] C1147;
wire A1147;
wire signed [6:0] C1207;
wire A1207;
wire signed [6:0] C1217;
wire A1217;
wire signed [6:0] C1227;
wire A1227;
wire signed [6:0] C1237;
wire A1237;
wire signed [6:0] C1247;
wire A1247;
wire signed [6:0] C1307;
wire A1307;
wire signed [6:0] C1317;
wire A1317;
wire signed [6:0] C1327;
wire A1327;
wire signed [6:0] C1337;
wire A1337;
wire signed [6:0] C1347;
wire A1347;
wire signed [6:0] C1407;
wire A1407;
wire signed [6:0] C1417;
wire A1417;
wire signed [6:0] C1427;
wire A1427;
wire signed [6:0] C1437;
wire A1437;
wire signed [6:0] C1447;
wire A1447;
wire signed [6:0] C1008;
wire A1008;
wire signed [6:0] C1018;
wire A1018;
wire signed [6:0] C1028;
wire A1028;
wire signed [6:0] C1038;
wire A1038;
wire signed [6:0] C1048;
wire A1048;
wire signed [6:0] C1108;
wire A1108;
wire signed [6:0] C1118;
wire A1118;
wire signed [6:0] C1128;
wire A1128;
wire signed [6:0] C1138;
wire A1138;
wire signed [6:0] C1148;
wire A1148;
wire signed [6:0] C1208;
wire A1208;
wire signed [6:0] C1218;
wire A1218;
wire signed [6:0] C1228;
wire A1228;
wire signed [6:0] C1238;
wire A1238;
wire signed [6:0] C1248;
wire A1248;
wire signed [6:0] C1308;
wire A1308;
wire signed [6:0] C1318;
wire A1318;
wire signed [6:0] C1328;
wire A1328;
wire signed [6:0] C1338;
wire A1338;
wire signed [6:0] C1348;
wire A1348;
wire signed [6:0] C1408;
wire A1408;
wire signed [6:0] C1418;
wire A1418;
wire signed [6:0] C1428;
wire A1428;
wire signed [6:0] C1438;
wire A1438;
wire signed [6:0] C1448;
wire A1448;
wire signed [6:0] C1009;
wire A1009;
wire signed [6:0] C1019;
wire A1019;
wire signed [6:0] C1029;
wire A1029;
wire signed [6:0] C1039;
wire A1039;
wire signed [6:0] C1049;
wire A1049;
wire signed [6:0] C1109;
wire A1109;
wire signed [6:0] C1119;
wire A1119;
wire signed [6:0] C1129;
wire A1129;
wire signed [6:0] C1139;
wire A1139;
wire signed [6:0] C1149;
wire A1149;
wire signed [6:0] C1209;
wire A1209;
wire signed [6:0] C1219;
wire A1219;
wire signed [6:0] C1229;
wire A1229;
wire signed [6:0] C1239;
wire A1239;
wire signed [6:0] C1249;
wire A1249;
wire signed [6:0] C1309;
wire A1309;
wire signed [6:0] C1319;
wire A1319;
wire signed [6:0] C1329;
wire A1329;
wire signed [6:0] C1339;
wire A1339;
wire signed [6:0] C1349;
wire A1349;
wire signed [6:0] C1409;
wire A1409;
wire signed [6:0] C1419;
wire A1419;
wire signed [6:0] C1429;
wire A1429;
wire signed [6:0] C1439;
wire A1439;
wire signed [6:0] C1449;
wire A1449;
wire signed [6:0] C100A;
wire A100A;
wire signed [6:0] C101A;
wire A101A;
wire signed [6:0] C102A;
wire A102A;
wire signed [6:0] C103A;
wire A103A;
wire signed [6:0] C104A;
wire A104A;
wire signed [6:0] C110A;
wire A110A;
wire signed [6:0] C111A;
wire A111A;
wire signed [6:0] C112A;
wire A112A;
wire signed [6:0] C113A;
wire A113A;
wire signed [6:0] C114A;
wire A114A;
wire signed [6:0] C120A;
wire A120A;
wire signed [6:0] C121A;
wire A121A;
wire signed [6:0] C122A;
wire A122A;
wire signed [6:0] C123A;
wire A123A;
wire signed [6:0] C124A;
wire A124A;
wire signed [6:0] C130A;
wire A130A;
wire signed [6:0] C131A;
wire A131A;
wire signed [6:0] C132A;
wire A132A;
wire signed [6:0] C133A;
wire A133A;
wire signed [6:0] C134A;
wire A134A;
wire signed [6:0] C140A;
wire A140A;
wire signed [6:0] C141A;
wire A141A;
wire signed [6:0] C142A;
wire A142A;
wire signed [6:0] C143A;
wire A143A;
wire signed [6:0] C144A;
wire A144A;
wire signed [6:0] C100B;
wire A100B;
wire signed [6:0] C101B;
wire A101B;
wire signed [6:0] C102B;
wire A102B;
wire signed [6:0] C103B;
wire A103B;
wire signed [6:0] C104B;
wire A104B;
wire signed [6:0] C110B;
wire A110B;
wire signed [6:0] C111B;
wire A111B;
wire signed [6:0] C112B;
wire A112B;
wire signed [6:0] C113B;
wire A113B;
wire signed [6:0] C114B;
wire A114B;
wire signed [6:0] C120B;
wire A120B;
wire signed [6:0] C121B;
wire A121B;
wire signed [6:0] C122B;
wire A122B;
wire signed [6:0] C123B;
wire A123B;
wire signed [6:0] C124B;
wire A124B;
wire signed [6:0] C130B;
wire A130B;
wire signed [6:0] C131B;
wire A131B;
wire signed [6:0] C132B;
wire A132B;
wire signed [6:0] C133B;
wire A133B;
wire signed [6:0] C134B;
wire A134B;
wire signed [6:0] C140B;
wire A140B;
wire signed [6:0] C141B;
wire A141B;
wire signed [6:0] C142B;
wire A142B;
wire signed [6:0] C143B;
wire A143B;
wire signed [6:0] C144B;
wire A144B;
wire signed [6:0] C100C;
wire A100C;
wire signed [6:0] C101C;
wire A101C;
wire signed [6:0] C102C;
wire A102C;
wire signed [6:0] C103C;
wire A103C;
wire signed [6:0] C104C;
wire A104C;
wire signed [6:0] C110C;
wire A110C;
wire signed [6:0] C111C;
wire A111C;
wire signed [6:0] C112C;
wire A112C;
wire signed [6:0] C113C;
wire A113C;
wire signed [6:0] C114C;
wire A114C;
wire signed [6:0] C120C;
wire A120C;
wire signed [6:0] C121C;
wire A121C;
wire signed [6:0] C122C;
wire A122C;
wire signed [6:0] C123C;
wire A123C;
wire signed [6:0] C124C;
wire A124C;
wire signed [6:0] C130C;
wire A130C;
wire signed [6:0] C131C;
wire A131C;
wire signed [6:0] C132C;
wire A132C;
wire signed [6:0] C133C;
wire A133C;
wire signed [6:0] C134C;
wire A134C;
wire signed [6:0] C140C;
wire A140C;
wire signed [6:0] C141C;
wire A141C;
wire signed [6:0] C142C;
wire A142C;
wire signed [6:0] C143C;
wire A143C;
wire signed [6:0] C144C;
wire A144C;
wire signed [6:0] C100D;
wire A100D;
wire signed [6:0] C101D;
wire A101D;
wire signed [6:0] C102D;
wire A102D;
wire signed [6:0] C103D;
wire A103D;
wire signed [6:0] C104D;
wire A104D;
wire signed [6:0] C110D;
wire A110D;
wire signed [6:0] C111D;
wire A111D;
wire signed [6:0] C112D;
wire A112D;
wire signed [6:0] C113D;
wire A113D;
wire signed [6:0] C114D;
wire A114D;
wire signed [6:0] C120D;
wire A120D;
wire signed [6:0] C121D;
wire A121D;
wire signed [6:0] C122D;
wire A122D;
wire signed [6:0] C123D;
wire A123D;
wire signed [6:0] C124D;
wire A124D;
wire signed [6:0] C130D;
wire A130D;
wire signed [6:0] C131D;
wire A131D;
wire signed [6:0] C132D;
wire A132D;
wire signed [6:0] C133D;
wire A133D;
wire signed [6:0] C134D;
wire A134D;
wire signed [6:0] C140D;
wire A140D;
wire signed [6:0] C141D;
wire A141D;
wire signed [6:0] C142D;
wire A142D;
wire signed [6:0] C143D;
wire A143D;
wire signed [6:0] C144D;
wire A144D;
wire signed [6:0] C100E;
wire A100E;
wire signed [6:0] C101E;
wire A101E;
wire signed [6:0] C102E;
wire A102E;
wire signed [6:0] C103E;
wire A103E;
wire signed [6:0] C104E;
wire A104E;
wire signed [6:0] C110E;
wire A110E;
wire signed [6:0] C111E;
wire A111E;
wire signed [6:0] C112E;
wire A112E;
wire signed [6:0] C113E;
wire A113E;
wire signed [6:0] C114E;
wire A114E;
wire signed [6:0] C120E;
wire A120E;
wire signed [6:0] C121E;
wire A121E;
wire signed [6:0] C122E;
wire A122E;
wire signed [6:0] C123E;
wire A123E;
wire signed [6:0] C124E;
wire A124E;
wire signed [6:0] C130E;
wire A130E;
wire signed [6:0] C131E;
wire A131E;
wire signed [6:0] C132E;
wire A132E;
wire signed [6:0] C133E;
wire A133E;
wire signed [6:0] C134E;
wire A134E;
wire signed [6:0] C140E;
wire A140E;
wire signed [6:0] C141E;
wire A141E;
wire signed [6:0] C142E;
wire A142E;
wire signed [6:0] C143E;
wire A143E;
wire signed [6:0] C144E;
wire A144E;
wire signed [6:0] C100F;
wire A100F;
wire signed [6:0] C101F;
wire A101F;
wire signed [6:0] C102F;
wire A102F;
wire signed [6:0] C103F;
wire A103F;
wire signed [6:0] C104F;
wire A104F;
wire signed [6:0] C110F;
wire A110F;
wire signed [6:0] C111F;
wire A111F;
wire signed [6:0] C112F;
wire A112F;
wire signed [6:0] C113F;
wire A113F;
wire signed [6:0] C114F;
wire A114F;
wire signed [6:0] C120F;
wire A120F;
wire signed [6:0] C121F;
wire A121F;
wire signed [6:0] C122F;
wire A122F;
wire signed [6:0] C123F;
wire A123F;
wire signed [6:0] C124F;
wire A124F;
wire signed [6:0] C130F;
wire A130F;
wire signed [6:0] C131F;
wire A131F;
wire signed [6:0] C132F;
wire A132F;
wire signed [6:0] C133F;
wire A133F;
wire signed [6:0] C134F;
wire A134F;
wire signed [6:0] C140F;
wire A140F;
wire signed [6:0] C141F;
wire A141F;
wire signed [6:0] C142F;
wire A142F;
wire signed [6:0] C143F;
wire A143F;
wire signed [6:0] C144F;
wire A144F;
DFF_save_fm DFF_W81(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10000));
DFF_save_fm DFF_W82(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10010));
DFF_save_fm DFF_W83(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10020));
DFF_save_fm DFF_W84(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10100));
DFF_save_fm DFF_W85(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10110));
DFF_save_fm DFF_W86(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10120));
DFF_save_fm DFF_W87(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10200));
DFF_save_fm DFF_W88(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10210));
DFF_save_fm DFF_W89(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10220));
DFF_save_fm DFF_W90(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10001));
DFF_save_fm DFF_W91(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10011));
DFF_save_fm DFF_W92(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10021));
DFF_save_fm DFF_W93(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10101));
DFF_save_fm DFF_W94(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10111));
DFF_save_fm DFF_W95(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10121));
DFF_save_fm DFF_W96(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10201));
DFF_save_fm DFF_W97(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10211));
DFF_save_fm DFF_W98(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10221));
DFF_save_fm DFF_W99(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10002));
DFF_save_fm DFF_W100(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10012));
DFF_save_fm DFF_W101(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10022));
DFF_save_fm DFF_W102(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10102));
DFF_save_fm DFF_W103(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10112));
DFF_save_fm DFF_W104(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10122));
DFF_save_fm DFF_W105(.clk(clk),.rstn(rstn),.reset_value(0),.q(W10202));
DFF_save_fm DFF_W106(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10212));
DFF_save_fm DFF_W107(.clk(clk),.rstn(rstn),.reset_value(1),.q(W10222));
DFF_save_fm DFF_W108(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11000));
DFF_save_fm DFF_W109(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11010));
DFF_save_fm DFF_W110(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11020));
DFF_save_fm DFF_W111(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11100));
DFF_save_fm DFF_W112(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11110));
DFF_save_fm DFF_W113(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11120));
DFF_save_fm DFF_W114(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11200));
DFF_save_fm DFF_W115(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11210));
DFF_save_fm DFF_W116(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11220));
DFF_save_fm DFF_W117(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11001));
DFF_save_fm DFF_W118(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11011));
DFF_save_fm DFF_W119(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11021));
DFF_save_fm DFF_W120(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11101));
DFF_save_fm DFF_W121(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11111));
DFF_save_fm DFF_W122(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11121));
DFF_save_fm DFF_W123(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11201));
DFF_save_fm DFF_W124(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11211));
DFF_save_fm DFF_W125(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11221));
DFF_save_fm DFF_W126(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11002));
DFF_save_fm DFF_W127(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11012));
DFF_save_fm DFF_W128(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11022));
DFF_save_fm DFF_W129(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11102));
DFF_save_fm DFF_W130(.clk(clk),.rstn(rstn),.reset_value(0),.q(W11112));
DFF_save_fm DFF_W131(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11122));
DFF_save_fm DFF_W132(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11202));
DFF_save_fm DFF_W133(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11212));
DFF_save_fm DFF_W134(.clk(clk),.rstn(rstn),.reset_value(1),.q(W11222));
DFF_save_fm DFF_W135(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12000));
DFF_save_fm DFF_W136(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12010));
DFF_save_fm DFF_W137(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12020));
DFF_save_fm DFF_W138(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12100));
DFF_save_fm DFF_W139(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12110));
DFF_save_fm DFF_W140(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12120));
DFF_save_fm DFF_W141(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12200));
DFF_save_fm DFF_W142(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12210));
DFF_save_fm DFF_W143(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12220));
DFF_save_fm DFF_W144(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12001));
DFF_save_fm DFF_W145(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12011));
DFF_save_fm DFF_W146(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12021));
DFF_save_fm DFF_W147(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12101));
DFF_save_fm DFF_W148(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12111));
DFF_save_fm DFF_W149(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12121));
DFF_save_fm DFF_W150(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12201));
DFF_save_fm DFF_W151(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12211));
DFF_save_fm DFF_W152(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12221));
DFF_save_fm DFF_W153(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12002));
DFF_save_fm DFF_W154(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12012));
DFF_save_fm DFF_W155(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12022));
DFF_save_fm DFF_W156(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12102));
DFF_save_fm DFF_W157(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12112));
DFF_save_fm DFF_W158(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12122));
DFF_save_fm DFF_W159(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12202));
DFF_save_fm DFF_W160(.clk(clk),.rstn(rstn),.reset_value(0),.q(W12212));
DFF_save_fm DFF_W161(.clk(clk),.rstn(rstn),.reset_value(1),.q(W12222));
DFF_save_fm DFF_W162(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13000));
DFF_save_fm DFF_W163(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13010));
DFF_save_fm DFF_W164(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13020));
DFF_save_fm DFF_W165(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13100));
DFF_save_fm DFF_W166(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13110));
DFF_save_fm DFF_W167(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13120));
DFF_save_fm DFF_W168(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13200));
DFF_save_fm DFF_W169(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13210));
DFF_save_fm DFF_W170(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13220));
DFF_save_fm DFF_W171(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13001));
DFF_save_fm DFF_W172(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13011));
DFF_save_fm DFF_W173(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13021));
DFF_save_fm DFF_W174(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13101));
DFF_save_fm DFF_W175(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13111));
DFF_save_fm DFF_W176(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13121));
DFF_save_fm DFF_W177(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13201));
DFF_save_fm DFF_W178(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13211));
DFF_save_fm DFF_W179(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13221));
DFF_save_fm DFF_W180(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13002));
DFF_save_fm DFF_W181(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13012));
DFF_save_fm DFF_W182(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13022));
DFF_save_fm DFF_W183(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13102));
DFF_save_fm DFF_W184(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13112));
DFF_save_fm DFF_W185(.clk(clk),.rstn(rstn),.reset_value(1),.q(W13122));
DFF_save_fm DFF_W186(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13202));
DFF_save_fm DFF_W187(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13212));
DFF_save_fm DFF_W188(.clk(clk),.rstn(rstn),.reset_value(0),.q(W13222));
DFF_save_fm DFF_W189(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14000));
DFF_save_fm DFF_W190(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14010));
DFF_save_fm DFF_W191(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14020));
DFF_save_fm DFF_W192(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14100));
DFF_save_fm DFF_W193(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14110));
DFF_save_fm DFF_W194(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14120));
DFF_save_fm DFF_W195(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14200));
DFF_save_fm DFF_W196(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14210));
DFF_save_fm DFF_W197(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14220));
DFF_save_fm DFF_W198(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14001));
DFF_save_fm DFF_W199(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14011));
DFF_save_fm DFF_W200(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14021));
DFF_save_fm DFF_W201(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14101));
DFF_save_fm DFF_W202(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14111));
DFF_save_fm DFF_W203(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14121));
DFF_save_fm DFF_W204(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14201));
DFF_save_fm DFF_W205(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14211));
DFF_save_fm DFF_W206(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14221));
DFF_save_fm DFF_W207(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14002));
DFF_save_fm DFF_W208(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14012));
DFF_save_fm DFF_W209(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14022));
DFF_save_fm DFF_W210(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14102));
DFF_save_fm DFF_W211(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14112));
DFF_save_fm DFF_W212(.clk(clk),.rstn(rstn),.reset_value(0),.q(W14122));
DFF_save_fm DFF_W213(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14202));
DFF_save_fm DFF_W214(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14212));
DFF_save_fm DFF_W215(.clk(clk),.rstn(rstn),.reset_value(1),.q(W14222));
DFF_save_fm DFF_W216(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15000));
DFF_save_fm DFF_W217(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15010));
DFF_save_fm DFF_W218(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15020));
DFF_save_fm DFF_W219(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15100));
DFF_save_fm DFF_W220(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15110));
DFF_save_fm DFF_W221(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15120));
DFF_save_fm DFF_W222(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15200));
DFF_save_fm DFF_W223(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15210));
DFF_save_fm DFF_W224(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15220));
DFF_save_fm DFF_W225(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15001));
DFF_save_fm DFF_W226(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15011));
DFF_save_fm DFF_W227(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15021));
DFF_save_fm DFF_W228(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15101));
DFF_save_fm DFF_W229(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15111));
DFF_save_fm DFF_W230(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15121));
DFF_save_fm DFF_W231(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15201));
DFF_save_fm DFF_W232(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15211));
DFF_save_fm DFF_W233(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15221));
DFF_save_fm DFF_W234(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15002));
DFF_save_fm DFF_W235(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15012));
DFF_save_fm DFF_W236(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15022));
DFF_save_fm DFF_W237(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15102));
DFF_save_fm DFF_W238(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15112));
DFF_save_fm DFF_W239(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15122));
DFF_save_fm DFF_W240(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15202));
DFF_save_fm DFF_W241(.clk(clk),.rstn(rstn),.reset_value(0),.q(W15212));
DFF_save_fm DFF_W242(.clk(clk),.rstn(rstn),.reset_value(1),.q(W15222));
DFF_save_fm DFF_W243(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16000));
DFF_save_fm DFF_W244(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16010));
DFF_save_fm DFF_W245(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16020));
DFF_save_fm DFF_W246(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16100));
DFF_save_fm DFF_W247(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16110));
DFF_save_fm DFF_W248(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16120));
DFF_save_fm DFF_W249(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16200));
DFF_save_fm DFF_W250(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16210));
DFF_save_fm DFF_W251(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16220));
DFF_save_fm DFF_W252(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16001));
DFF_save_fm DFF_W253(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16011));
DFF_save_fm DFF_W254(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16021));
DFF_save_fm DFF_W255(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16101));
DFF_save_fm DFF_W256(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16111));
DFF_save_fm DFF_W257(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16121));
DFF_save_fm DFF_W258(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16201));
DFF_save_fm DFF_W259(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16211));
DFF_save_fm DFF_W260(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16221));
DFF_save_fm DFF_W261(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16002));
DFF_save_fm DFF_W262(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16012));
DFF_save_fm DFF_W263(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16022));
DFF_save_fm DFF_W264(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16102));
DFF_save_fm DFF_W265(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16112));
DFF_save_fm DFF_W266(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16122));
DFF_save_fm DFF_W267(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16202));
DFF_save_fm DFF_W268(.clk(clk),.rstn(rstn),.reset_value(1),.q(W16212));
DFF_save_fm DFF_W269(.clk(clk),.rstn(rstn),.reset_value(0),.q(W16222));
DFF_save_fm DFF_W270(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17000));
DFF_save_fm DFF_W271(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17010));
DFF_save_fm DFF_W272(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17020));
DFF_save_fm DFF_W273(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17100));
DFF_save_fm DFF_W274(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17110));
DFF_save_fm DFF_W275(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17120));
DFF_save_fm DFF_W276(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17200));
DFF_save_fm DFF_W277(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17210));
DFF_save_fm DFF_W278(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17220));
DFF_save_fm DFF_W279(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17001));
DFF_save_fm DFF_W280(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17011));
DFF_save_fm DFF_W281(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17021));
DFF_save_fm DFF_W282(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17101));
DFF_save_fm DFF_W283(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17111));
DFF_save_fm DFF_W284(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17121));
DFF_save_fm DFF_W285(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17201));
DFF_save_fm DFF_W286(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17211));
DFF_save_fm DFF_W287(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17221));
DFF_save_fm DFF_W288(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17002));
DFF_save_fm DFF_W289(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17012));
DFF_save_fm DFF_W290(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17022));
DFF_save_fm DFF_W291(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17102));
DFF_save_fm DFF_W292(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17112));
DFF_save_fm DFF_W293(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17122));
DFF_save_fm DFF_W294(.clk(clk),.rstn(rstn),.reset_value(1),.q(W17202));
DFF_save_fm DFF_W295(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17212));
DFF_save_fm DFF_W296(.clk(clk),.rstn(rstn),.reset_value(0),.q(W17222));
DFF_save_fm DFF_W297(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18000));
DFF_save_fm DFF_W298(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18010));
DFF_save_fm DFF_W299(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18020));
DFF_save_fm DFF_W300(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18100));
DFF_save_fm DFF_W301(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18110));
DFF_save_fm DFF_W302(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18120));
DFF_save_fm DFF_W303(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18200));
DFF_save_fm DFF_W304(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18210));
DFF_save_fm DFF_W305(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18220));
DFF_save_fm DFF_W306(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18001));
DFF_save_fm DFF_W307(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18011));
DFF_save_fm DFF_W308(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18021));
DFF_save_fm DFF_W309(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18101));
DFF_save_fm DFF_W310(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18111));
DFF_save_fm DFF_W311(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18121));
DFF_save_fm DFF_W312(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18201));
DFF_save_fm DFF_W313(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18211));
DFF_save_fm DFF_W314(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18221));
DFF_save_fm DFF_W315(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18002));
DFF_save_fm DFF_W316(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18012));
DFF_save_fm DFF_W317(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18022));
DFF_save_fm DFF_W318(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18102));
DFF_save_fm DFF_W319(.clk(clk),.rstn(rstn),.reset_value(1),.q(W18112));
DFF_save_fm DFF_W320(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18122));
DFF_save_fm DFF_W321(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18202));
DFF_save_fm DFF_W322(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18212));
DFF_save_fm DFF_W323(.clk(clk),.rstn(rstn),.reset_value(0),.q(W18222));
DFF_save_fm DFF_W324(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19000));
DFF_save_fm DFF_W325(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19010));
DFF_save_fm DFF_W326(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19020));
DFF_save_fm DFF_W327(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19100));
DFF_save_fm DFF_W328(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19110));
DFF_save_fm DFF_W329(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19120));
DFF_save_fm DFF_W330(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19200));
DFF_save_fm DFF_W331(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19210));
DFF_save_fm DFF_W332(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19220));
DFF_save_fm DFF_W333(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19001));
DFF_save_fm DFF_W334(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19011));
DFF_save_fm DFF_W335(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19021));
DFF_save_fm DFF_W336(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19101));
DFF_save_fm DFF_W337(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19111));
DFF_save_fm DFF_W338(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19121));
DFF_save_fm DFF_W339(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19201));
DFF_save_fm DFF_W340(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19211));
DFF_save_fm DFF_W341(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19221));
DFF_save_fm DFF_W342(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19002));
DFF_save_fm DFF_W343(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19012));
DFF_save_fm DFF_W344(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19022));
DFF_save_fm DFF_W345(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19102));
DFF_save_fm DFF_W346(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19112));
DFF_save_fm DFF_W347(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19122));
DFF_save_fm DFF_W348(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19202));
DFF_save_fm DFF_W349(.clk(clk),.rstn(rstn),.reset_value(0),.q(W19212));
DFF_save_fm DFF_W350(.clk(clk),.rstn(rstn),.reset_value(1),.q(W19222));
DFF_save_fm DFF_W351(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A000));
DFF_save_fm DFF_W352(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A010));
DFF_save_fm DFF_W353(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A020));
DFF_save_fm DFF_W354(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A100));
DFF_save_fm DFF_W355(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A110));
DFF_save_fm DFF_W356(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A120));
DFF_save_fm DFF_W357(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A200));
DFF_save_fm DFF_W358(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A210));
DFF_save_fm DFF_W359(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A220));
DFF_save_fm DFF_W360(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A001));
DFF_save_fm DFF_W361(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A011));
DFF_save_fm DFF_W362(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A021));
DFF_save_fm DFF_W363(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A101));
DFF_save_fm DFF_W364(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A111));
DFF_save_fm DFF_W365(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A121));
DFF_save_fm DFF_W366(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A201));
DFF_save_fm DFF_W367(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A211));
DFF_save_fm DFF_W368(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A221));
DFF_save_fm DFF_W369(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A002));
DFF_save_fm DFF_W370(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A012));
DFF_save_fm DFF_W371(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A022));
DFF_save_fm DFF_W372(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A102));
DFF_save_fm DFF_W373(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A112));
DFF_save_fm DFF_W374(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A122));
DFF_save_fm DFF_W375(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A202));
DFF_save_fm DFF_W376(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1A212));
DFF_save_fm DFF_W377(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1A222));
DFF_save_fm DFF_W378(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B000));
DFF_save_fm DFF_W379(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B010));
DFF_save_fm DFF_W380(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B020));
DFF_save_fm DFF_W381(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B100));
DFF_save_fm DFF_W382(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B110));
DFF_save_fm DFF_W383(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B120));
DFF_save_fm DFF_W384(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B200));
DFF_save_fm DFF_W385(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B210));
DFF_save_fm DFF_W386(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B220));
DFF_save_fm DFF_W387(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B001));
DFF_save_fm DFF_W388(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B011));
DFF_save_fm DFF_W389(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B021));
DFF_save_fm DFF_W390(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B101));
DFF_save_fm DFF_W391(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B111));
DFF_save_fm DFF_W392(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B121));
DFF_save_fm DFF_W393(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B201));
DFF_save_fm DFF_W394(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B211));
DFF_save_fm DFF_W395(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B221));
DFF_save_fm DFF_W396(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B002));
DFF_save_fm DFF_W397(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B012));
DFF_save_fm DFF_W398(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B022));
DFF_save_fm DFF_W399(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B102));
DFF_save_fm DFF_W400(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B112));
DFF_save_fm DFF_W401(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B122));
DFF_save_fm DFF_W402(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1B202));
DFF_save_fm DFF_W403(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B212));
DFF_save_fm DFF_W404(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1B222));
DFF_save_fm DFF_W405(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C000));
DFF_save_fm DFF_W406(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C010));
DFF_save_fm DFF_W407(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C020));
DFF_save_fm DFF_W408(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C100));
DFF_save_fm DFF_W409(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C110));
DFF_save_fm DFF_W410(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C120));
DFF_save_fm DFF_W411(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C200));
DFF_save_fm DFF_W412(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C210));
DFF_save_fm DFF_W413(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C220));
DFF_save_fm DFF_W414(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C001));
DFF_save_fm DFF_W415(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C011));
DFF_save_fm DFF_W416(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C021));
DFF_save_fm DFF_W417(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C101));
DFF_save_fm DFF_W418(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C111));
DFF_save_fm DFF_W419(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C121));
DFF_save_fm DFF_W420(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C201));
DFF_save_fm DFF_W421(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C211));
DFF_save_fm DFF_W422(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C221));
DFF_save_fm DFF_W423(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C002));
DFF_save_fm DFF_W424(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C012));
DFF_save_fm DFF_W425(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C022));
DFF_save_fm DFF_W426(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C102));
DFF_save_fm DFF_W427(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C112));
DFF_save_fm DFF_W428(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1C122));
DFF_save_fm DFF_W429(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C202));
DFF_save_fm DFF_W430(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C212));
DFF_save_fm DFF_W431(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1C222));
DFF_save_fm DFF_W432(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D000));
DFF_save_fm DFF_W433(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D010));
DFF_save_fm DFF_W434(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D020));
DFF_save_fm DFF_W435(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D100));
DFF_save_fm DFF_W436(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D110));
DFF_save_fm DFF_W437(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D120));
DFF_save_fm DFF_W438(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D200));
DFF_save_fm DFF_W439(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D210));
DFF_save_fm DFF_W440(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D220));
DFF_save_fm DFF_W441(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D001));
DFF_save_fm DFF_W442(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D011));
DFF_save_fm DFF_W443(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D021));
DFF_save_fm DFF_W444(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D101));
DFF_save_fm DFF_W445(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D111));
DFF_save_fm DFF_W446(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D121));
DFF_save_fm DFF_W447(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D201));
DFF_save_fm DFF_W448(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D211));
DFF_save_fm DFF_W449(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D221));
DFF_save_fm DFF_W450(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D002));
DFF_save_fm DFF_W451(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D012));
DFF_save_fm DFF_W452(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D022));
DFF_save_fm DFF_W453(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D102));
DFF_save_fm DFF_W454(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D112));
DFF_save_fm DFF_W455(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D122));
DFF_save_fm DFF_W456(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D202));
DFF_save_fm DFF_W457(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1D212));
DFF_save_fm DFF_W458(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1D222));
DFF_save_fm DFF_W459(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E000));
DFF_save_fm DFF_W460(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E010));
DFF_save_fm DFF_W461(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E020));
DFF_save_fm DFF_W462(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E100));
DFF_save_fm DFF_W463(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E110));
DFF_save_fm DFF_W464(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E120));
DFF_save_fm DFF_W465(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E200));
DFF_save_fm DFF_W466(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E210));
DFF_save_fm DFF_W467(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E220));
DFF_save_fm DFF_W468(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E001));
DFF_save_fm DFF_W469(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E011));
DFF_save_fm DFF_W470(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E021));
DFF_save_fm DFF_W471(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E101));
DFF_save_fm DFF_W472(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E111));
DFF_save_fm DFF_W473(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E121));
DFF_save_fm DFF_W474(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E201));
DFF_save_fm DFF_W475(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E211));
DFF_save_fm DFF_W476(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E221));
DFF_save_fm DFF_W477(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E002));
DFF_save_fm DFF_W478(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E012));
DFF_save_fm DFF_W479(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E022));
DFF_save_fm DFF_W480(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E102));
DFF_save_fm DFF_W481(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E112));
DFF_save_fm DFF_W482(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E122));
DFF_save_fm DFF_W483(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E202));
DFF_save_fm DFF_W484(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1E212));
DFF_save_fm DFF_W485(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1E222));
DFF_save_fm DFF_W486(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F000));
DFF_save_fm DFF_W487(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F010));
DFF_save_fm DFF_W488(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F020));
DFF_save_fm DFF_W489(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F100));
DFF_save_fm DFF_W490(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F110));
DFF_save_fm DFF_W491(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F120));
DFF_save_fm DFF_W492(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F200));
DFF_save_fm DFF_W493(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F210));
DFF_save_fm DFF_W494(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F220));
DFF_save_fm DFF_W495(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F001));
DFF_save_fm DFF_W496(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F011));
DFF_save_fm DFF_W497(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F021));
DFF_save_fm DFF_W498(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F101));
DFF_save_fm DFF_W499(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F111));
DFF_save_fm DFF_W500(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F121));
DFF_save_fm DFF_W501(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F201));
DFF_save_fm DFF_W502(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F211));
DFF_save_fm DFF_W503(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F221));
DFF_save_fm DFF_W504(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F002));
DFF_save_fm DFF_W505(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F012));
DFF_save_fm DFF_W506(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F022));
DFF_save_fm DFF_W507(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F102));
DFF_save_fm DFF_W508(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F112));
DFF_save_fm DFF_W509(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F122));
DFF_save_fm DFF_W510(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F202));
DFF_save_fm DFF_W511(.clk(clk),.rstn(rstn),.reset_value(1),.q(W1F212));
DFF_save_fm DFF_W512(.clk(clk),.rstn(rstn),.reset_value(0),.q(W1F222));
ninexnine_unit ninexnine_unit_1764(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10000)
);

ninexnine_unit ninexnine_unit_1765(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11000)
);

ninexnine_unit ninexnine_unit_1766(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12000)
);

assign C1000=c10000+c11000+c12000;
assign A1000=(C1000>=0)?1:0;

assign P2000=A1000;

ninexnine_unit ninexnine_unit_1767(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10010)
);

ninexnine_unit ninexnine_unit_1768(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11010)
);

ninexnine_unit ninexnine_unit_1769(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12010)
);

assign C1010=c10010+c11010+c12010;
assign A1010=(C1010>=0)?1:0;

assign P2010=A1010;

ninexnine_unit ninexnine_unit_1770(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10020)
);

ninexnine_unit ninexnine_unit_1771(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11020)
);

ninexnine_unit ninexnine_unit_1772(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12020)
);

assign C1020=c10020+c11020+c12020;
assign A1020=(C1020>=0)?1:0;

assign P2020=A1020;

ninexnine_unit ninexnine_unit_1773(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10030)
);

ninexnine_unit ninexnine_unit_1774(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11030)
);

ninexnine_unit ninexnine_unit_1775(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12030)
);

assign C1030=c10030+c11030+c12030;
assign A1030=(C1030>=0)?1:0;

assign P2030=A1030;

ninexnine_unit ninexnine_unit_1776(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10040)
);

ninexnine_unit ninexnine_unit_1777(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11040)
);

ninexnine_unit ninexnine_unit_1778(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12040)
);

assign C1040=c10040+c11040+c12040;
assign A1040=(C1040>=0)?1:0;

assign P2040=A1040;

ninexnine_unit ninexnine_unit_1779(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10100)
);

ninexnine_unit ninexnine_unit_1780(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11100)
);

ninexnine_unit ninexnine_unit_1781(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12100)
);

assign C1100=c10100+c11100+c12100;
assign A1100=(C1100>=0)?1:0;

assign P2100=A1100;

ninexnine_unit ninexnine_unit_1782(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10110)
);

ninexnine_unit ninexnine_unit_1783(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11110)
);

ninexnine_unit ninexnine_unit_1784(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12110)
);

assign C1110=c10110+c11110+c12110;
assign A1110=(C1110>=0)?1:0;

assign P2110=A1110;

ninexnine_unit ninexnine_unit_1785(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10120)
);

ninexnine_unit ninexnine_unit_1786(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11120)
);

ninexnine_unit ninexnine_unit_1787(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12120)
);

assign C1120=c10120+c11120+c12120;
assign A1120=(C1120>=0)?1:0;

assign P2120=A1120;

ninexnine_unit ninexnine_unit_1788(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10130)
);

ninexnine_unit ninexnine_unit_1789(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11130)
);

ninexnine_unit ninexnine_unit_1790(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12130)
);

assign C1130=c10130+c11130+c12130;
assign A1130=(C1130>=0)?1:0;

assign P2130=A1130;

ninexnine_unit ninexnine_unit_1791(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10140)
);

ninexnine_unit ninexnine_unit_1792(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11140)
);

ninexnine_unit ninexnine_unit_1793(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12140)
);

assign C1140=c10140+c11140+c12140;
assign A1140=(C1140>=0)?1:0;

assign P2140=A1140;

ninexnine_unit ninexnine_unit_1794(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10200)
);

ninexnine_unit ninexnine_unit_1795(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11200)
);

ninexnine_unit ninexnine_unit_1796(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12200)
);

assign C1200=c10200+c11200+c12200;
assign A1200=(C1200>=0)?1:0;

assign P2200=A1200;

ninexnine_unit ninexnine_unit_1797(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10210)
);

ninexnine_unit ninexnine_unit_1798(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11210)
);

ninexnine_unit ninexnine_unit_1799(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12210)
);

assign C1210=c10210+c11210+c12210;
assign A1210=(C1210>=0)?1:0;

assign P2210=A1210;

ninexnine_unit ninexnine_unit_1800(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10220)
);

ninexnine_unit ninexnine_unit_1801(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11220)
);

ninexnine_unit ninexnine_unit_1802(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12220)
);

assign C1220=c10220+c11220+c12220;
assign A1220=(C1220>=0)?1:0;

assign P2220=A1220;

ninexnine_unit ninexnine_unit_1803(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10230)
);

ninexnine_unit ninexnine_unit_1804(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11230)
);

ninexnine_unit ninexnine_unit_1805(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12230)
);

assign C1230=c10230+c11230+c12230;
assign A1230=(C1230>=0)?1:0;

assign P2230=A1230;

ninexnine_unit ninexnine_unit_1806(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10240)
);

ninexnine_unit ninexnine_unit_1807(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11240)
);

ninexnine_unit ninexnine_unit_1808(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12240)
);

assign C1240=c10240+c11240+c12240;
assign A1240=(C1240>=0)?1:0;

assign P2240=A1240;

ninexnine_unit ninexnine_unit_1809(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10300)
);

ninexnine_unit ninexnine_unit_1810(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11300)
);

ninexnine_unit ninexnine_unit_1811(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12300)
);

assign C1300=c10300+c11300+c12300;
assign A1300=(C1300>=0)?1:0;

assign P2300=A1300;

ninexnine_unit ninexnine_unit_1812(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10310)
);

ninexnine_unit ninexnine_unit_1813(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11310)
);

ninexnine_unit ninexnine_unit_1814(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12310)
);

assign C1310=c10310+c11310+c12310;
assign A1310=(C1310>=0)?1:0;

assign P2310=A1310;

ninexnine_unit ninexnine_unit_1815(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10320)
);

ninexnine_unit ninexnine_unit_1816(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11320)
);

ninexnine_unit ninexnine_unit_1817(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12320)
);

assign C1320=c10320+c11320+c12320;
assign A1320=(C1320>=0)?1:0;

assign P2320=A1320;

ninexnine_unit ninexnine_unit_1818(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10330)
);

ninexnine_unit ninexnine_unit_1819(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11330)
);

ninexnine_unit ninexnine_unit_1820(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12330)
);

assign C1330=c10330+c11330+c12330;
assign A1330=(C1330>=0)?1:0;

assign P2330=A1330;

ninexnine_unit ninexnine_unit_1821(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10340)
);

ninexnine_unit ninexnine_unit_1822(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11340)
);

ninexnine_unit ninexnine_unit_1823(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12340)
);

assign C1340=c10340+c11340+c12340;
assign A1340=(C1340>=0)?1:0;

assign P2340=A1340;

ninexnine_unit ninexnine_unit_1824(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10400)
);

ninexnine_unit ninexnine_unit_1825(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11400)
);

ninexnine_unit ninexnine_unit_1826(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12400)
);

assign C1400=c10400+c11400+c12400;
assign A1400=(C1400>=0)?1:0;

assign P2400=A1400;

ninexnine_unit ninexnine_unit_1827(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10410)
);

ninexnine_unit ninexnine_unit_1828(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11410)
);

ninexnine_unit ninexnine_unit_1829(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12410)
);

assign C1410=c10410+c11410+c12410;
assign A1410=(C1410>=0)?1:0;

assign P2410=A1410;

ninexnine_unit ninexnine_unit_1830(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10420)
);

ninexnine_unit ninexnine_unit_1831(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11420)
);

ninexnine_unit ninexnine_unit_1832(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12420)
);

assign C1420=c10420+c11420+c12420;
assign A1420=(C1420>=0)?1:0;

assign P2420=A1420;

ninexnine_unit ninexnine_unit_1833(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10430)
);

ninexnine_unit ninexnine_unit_1834(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11430)
);

ninexnine_unit ninexnine_unit_1835(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12430)
);

assign C1430=c10430+c11430+c12430;
assign A1430=(C1430>=0)?1:0;

assign P2430=A1430;

ninexnine_unit ninexnine_unit_1836(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W10000),
				.b1(W10010),
				.b2(W10020),
				.b3(W10100),
				.b4(W10110),
				.b5(W10120),
				.b6(W10200),
				.b7(W10210),
				.b8(W10220),
				.c(c10440)
);

ninexnine_unit ninexnine_unit_1837(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W10001),
				.b1(W10011),
				.b2(W10021),
				.b3(W10101),
				.b4(W10111),
				.b5(W10121),
				.b6(W10201),
				.b7(W10211),
				.b8(W10221),
				.c(c11440)
);

ninexnine_unit ninexnine_unit_1838(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W10002),
				.b1(W10012),
				.b2(W10022),
				.b3(W10102),
				.b4(W10112),
				.b5(W10122),
				.b6(W10202),
				.b7(W10212),
				.b8(W10222),
				.c(c12440)
);

assign C1440=c10440+c11440+c12440;
assign A1440=(C1440>=0)?1:0;

assign P2440=A1440;

ninexnine_unit ninexnine_unit_1839(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10001)
);

ninexnine_unit ninexnine_unit_1840(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11001)
);

ninexnine_unit ninexnine_unit_1841(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12001)
);

assign C1001=c10001+c11001+c12001;
assign A1001=(C1001>=0)?1:0;

assign P2001=A1001;

ninexnine_unit ninexnine_unit_1842(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10011)
);

ninexnine_unit ninexnine_unit_1843(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11011)
);

ninexnine_unit ninexnine_unit_1844(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12011)
);

assign C1011=c10011+c11011+c12011;
assign A1011=(C1011>=0)?1:0;

assign P2011=A1011;

ninexnine_unit ninexnine_unit_1845(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10021)
);

ninexnine_unit ninexnine_unit_1846(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11021)
);

ninexnine_unit ninexnine_unit_1847(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12021)
);

assign C1021=c10021+c11021+c12021;
assign A1021=(C1021>=0)?1:0;

assign P2021=A1021;

ninexnine_unit ninexnine_unit_1848(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10031)
);

ninexnine_unit ninexnine_unit_1849(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11031)
);

ninexnine_unit ninexnine_unit_1850(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12031)
);

assign C1031=c10031+c11031+c12031;
assign A1031=(C1031>=0)?1:0;

assign P2031=A1031;

ninexnine_unit ninexnine_unit_1851(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10041)
);

ninexnine_unit ninexnine_unit_1852(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11041)
);

ninexnine_unit ninexnine_unit_1853(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12041)
);

assign C1041=c10041+c11041+c12041;
assign A1041=(C1041>=0)?1:0;

assign P2041=A1041;

ninexnine_unit ninexnine_unit_1854(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10101)
);

ninexnine_unit ninexnine_unit_1855(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11101)
);

ninexnine_unit ninexnine_unit_1856(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12101)
);

assign C1101=c10101+c11101+c12101;
assign A1101=(C1101>=0)?1:0;

assign P2101=A1101;

ninexnine_unit ninexnine_unit_1857(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10111)
);

ninexnine_unit ninexnine_unit_1858(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11111)
);

ninexnine_unit ninexnine_unit_1859(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12111)
);

assign C1111=c10111+c11111+c12111;
assign A1111=(C1111>=0)?1:0;

assign P2111=A1111;

ninexnine_unit ninexnine_unit_1860(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10121)
);

ninexnine_unit ninexnine_unit_1861(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11121)
);

ninexnine_unit ninexnine_unit_1862(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12121)
);

assign C1121=c10121+c11121+c12121;
assign A1121=(C1121>=0)?1:0;

assign P2121=A1121;

ninexnine_unit ninexnine_unit_1863(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10131)
);

ninexnine_unit ninexnine_unit_1864(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11131)
);

ninexnine_unit ninexnine_unit_1865(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12131)
);

assign C1131=c10131+c11131+c12131;
assign A1131=(C1131>=0)?1:0;

assign P2131=A1131;

ninexnine_unit ninexnine_unit_1866(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10141)
);

ninexnine_unit ninexnine_unit_1867(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11141)
);

ninexnine_unit ninexnine_unit_1868(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12141)
);

assign C1141=c10141+c11141+c12141;
assign A1141=(C1141>=0)?1:0;

assign P2141=A1141;

ninexnine_unit ninexnine_unit_1869(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10201)
);

ninexnine_unit ninexnine_unit_1870(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11201)
);

ninexnine_unit ninexnine_unit_1871(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12201)
);

assign C1201=c10201+c11201+c12201;
assign A1201=(C1201>=0)?1:0;

assign P2201=A1201;

ninexnine_unit ninexnine_unit_1872(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10211)
);

ninexnine_unit ninexnine_unit_1873(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11211)
);

ninexnine_unit ninexnine_unit_1874(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12211)
);

assign C1211=c10211+c11211+c12211;
assign A1211=(C1211>=0)?1:0;

assign P2211=A1211;

ninexnine_unit ninexnine_unit_1875(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10221)
);

ninexnine_unit ninexnine_unit_1876(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11221)
);

ninexnine_unit ninexnine_unit_1877(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12221)
);

assign C1221=c10221+c11221+c12221;
assign A1221=(C1221>=0)?1:0;

assign P2221=A1221;

ninexnine_unit ninexnine_unit_1878(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10231)
);

ninexnine_unit ninexnine_unit_1879(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11231)
);

ninexnine_unit ninexnine_unit_1880(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12231)
);

assign C1231=c10231+c11231+c12231;
assign A1231=(C1231>=0)?1:0;

assign P2231=A1231;

ninexnine_unit ninexnine_unit_1881(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10241)
);

ninexnine_unit ninexnine_unit_1882(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11241)
);

ninexnine_unit ninexnine_unit_1883(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12241)
);

assign C1241=c10241+c11241+c12241;
assign A1241=(C1241>=0)?1:0;

assign P2241=A1241;

ninexnine_unit ninexnine_unit_1884(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10301)
);

ninexnine_unit ninexnine_unit_1885(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11301)
);

ninexnine_unit ninexnine_unit_1886(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12301)
);

assign C1301=c10301+c11301+c12301;
assign A1301=(C1301>=0)?1:0;

assign P2301=A1301;

ninexnine_unit ninexnine_unit_1887(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10311)
);

ninexnine_unit ninexnine_unit_1888(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11311)
);

ninexnine_unit ninexnine_unit_1889(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12311)
);

assign C1311=c10311+c11311+c12311;
assign A1311=(C1311>=0)?1:0;

assign P2311=A1311;

ninexnine_unit ninexnine_unit_1890(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10321)
);

ninexnine_unit ninexnine_unit_1891(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11321)
);

ninexnine_unit ninexnine_unit_1892(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12321)
);

assign C1321=c10321+c11321+c12321;
assign A1321=(C1321>=0)?1:0;

assign P2321=A1321;

ninexnine_unit ninexnine_unit_1893(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10331)
);

ninexnine_unit ninexnine_unit_1894(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11331)
);

ninexnine_unit ninexnine_unit_1895(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12331)
);

assign C1331=c10331+c11331+c12331;
assign A1331=(C1331>=0)?1:0;

assign P2331=A1331;

ninexnine_unit ninexnine_unit_1896(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10341)
);

ninexnine_unit ninexnine_unit_1897(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11341)
);

ninexnine_unit ninexnine_unit_1898(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12341)
);

assign C1341=c10341+c11341+c12341;
assign A1341=(C1341>=0)?1:0;

assign P2341=A1341;

ninexnine_unit ninexnine_unit_1899(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10401)
);

ninexnine_unit ninexnine_unit_1900(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11401)
);

ninexnine_unit ninexnine_unit_1901(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12401)
);

assign C1401=c10401+c11401+c12401;
assign A1401=(C1401>=0)?1:0;

assign P2401=A1401;

ninexnine_unit ninexnine_unit_1902(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10411)
);

ninexnine_unit ninexnine_unit_1903(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11411)
);

ninexnine_unit ninexnine_unit_1904(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12411)
);

assign C1411=c10411+c11411+c12411;
assign A1411=(C1411>=0)?1:0;

assign P2411=A1411;

ninexnine_unit ninexnine_unit_1905(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10421)
);

ninexnine_unit ninexnine_unit_1906(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11421)
);

ninexnine_unit ninexnine_unit_1907(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12421)
);

assign C1421=c10421+c11421+c12421;
assign A1421=(C1421>=0)?1:0;

assign P2421=A1421;

ninexnine_unit ninexnine_unit_1908(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10431)
);

ninexnine_unit ninexnine_unit_1909(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11431)
);

ninexnine_unit ninexnine_unit_1910(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12431)
);

assign C1431=c10431+c11431+c12431;
assign A1431=(C1431>=0)?1:0;

assign P2431=A1431;

ninexnine_unit ninexnine_unit_1911(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W11000),
				.b1(W11010),
				.b2(W11020),
				.b3(W11100),
				.b4(W11110),
				.b5(W11120),
				.b6(W11200),
				.b7(W11210),
				.b8(W11220),
				.c(c10441)
);

ninexnine_unit ninexnine_unit_1912(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W11001),
				.b1(W11011),
				.b2(W11021),
				.b3(W11101),
				.b4(W11111),
				.b5(W11121),
				.b6(W11201),
				.b7(W11211),
				.b8(W11221),
				.c(c11441)
);

ninexnine_unit ninexnine_unit_1913(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W11002),
				.b1(W11012),
				.b2(W11022),
				.b3(W11102),
				.b4(W11112),
				.b5(W11122),
				.b6(W11202),
				.b7(W11212),
				.b8(W11222),
				.c(c12441)
);

assign C1441=c10441+c11441+c12441;
assign A1441=(C1441>=0)?1:0;

assign P2441=A1441;

ninexnine_unit ninexnine_unit_1914(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10002)
);

ninexnine_unit ninexnine_unit_1915(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11002)
);

ninexnine_unit ninexnine_unit_1916(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12002)
);

assign C1002=c10002+c11002+c12002;
assign A1002=(C1002>=0)?1:0;

assign P2002=A1002;

ninexnine_unit ninexnine_unit_1917(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10012)
);

ninexnine_unit ninexnine_unit_1918(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11012)
);

ninexnine_unit ninexnine_unit_1919(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12012)
);

assign C1012=c10012+c11012+c12012;
assign A1012=(C1012>=0)?1:0;

assign P2012=A1012;

ninexnine_unit ninexnine_unit_1920(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10022)
);

ninexnine_unit ninexnine_unit_1921(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11022)
);

ninexnine_unit ninexnine_unit_1922(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12022)
);

assign C1022=c10022+c11022+c12022;
assign A1022=(C1022>=0)?1:0;

assign P2022=A1022;

ninexnine_unit ninexnine_unit_1923(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10032)
);

ninexnine_unit ninexnine_unit_1924(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11032)
);

ninexnine_unit ninexnine_unit_1925(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12032)
);

assign C1032=c10032+c11032+c12032;
assign A1032=(C1032>=0)?1:0;

assign P2032=A1032;

ninexnine_unit ninexnine_unit_1926(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10042)
);

ninexnine_unit ninexnine_unit_1927(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11042)
);

ninexnine_unit ninexnine_unit_1928(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12042)
);

assign C1042=c10042+c11042+c12042;
assign A1042=(C1042>=0)?1:0;

assign P2042=A1042;

ninexnine_unit ninexnine_unit_1929(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10102)
);

ninexnine_unit ninexnine_unit_1930(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11102)
);

ninexnine_unit ninexnine_unit_1931(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12102)
);

assign C1102=c10102+c11102+c12102;
assign A1102=(C1102>=0)?1:0;

assign P2102=A1102;

ninexnine_unit ninexnine_unit_1932(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10112)
);

ninexnine_unit ninexnine_unit_1933(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11112)
);

ninexnine_unit ninexnine_unit_1934(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12112)
);

assign C1112=c10112+c11112+c12112;
assign A1112=(C1112>=0)?1:0;

assign P2112=A1112;

ninexnine_unit ninexnine_unit_1935(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10122)
);

ninexnine_unit ninexnine_unit_1936(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11122)
);

ninexnine_unit ninexnine_unit_1937(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12122)
);

assign C1122=c10122+c11122+c12122;
assign A1122=(C1122>=0)?1:0;

assign P2122=A1122;

ninexnine_unit ninexnine_unit_1938(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10132)
);

ninexnine_unit ninexnine_unit_1939(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11132)
);

ninexnine_unit ninexnine_unit_1940(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12132)
);

assign C1132=c10132+c11132+c12132;
assign A1132=(C1132>=0)?1:0;

assign P2132=A1132;

ninexnine_unit ninexnine_unit_1941(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10142)
);

ninexnine_unit ninexnine_unit_1942(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11142)
);

ninexnine_unit ninexnine_unit_1943(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12142)
);

assign C1142=c10142+c11142+c12142;
assign A1142=(C1142>=0)?1:0;

assign P2142=A1142;

ninexnine_unit ninexnine_unit_1944(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10202)
);

ninexnine_unit ninexnine_unit_1945(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11202)
);

ninexnine_unit ninexnine_unit_1946(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12202)
);

assign C1202=c10202+c11202+c12202;
assign A1202=(C1202>=0)?1:0;

assign P2202=A1202;

ninexnine_unit ninexnine_unit_1947(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10212)
);

ninexnine_unit ninexnine_unit_1948(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11212)
);

ninexnine_unit ninexnine_unit_1949(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12212)
);

assign C1212=c10212+c11212+c12212;
assign A1212=(C1212>=0)?1:0;

assign P2212=A1212;

ninexnine_unit ninexnine_unit_1950(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10222)
);

ninexnine_unit ninexnine_unit_1951(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11222)
);

ninexnine_unit ninexnine_unit_1952(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12222)
);

assign C1222=c10222+c11222+c12222;
assign A1222=(C1222>=0)?1:0;

assign P2222=A1222;

ninexnine_unit ninexnine_unit_1953(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10232)
);

ninexnine_unit ninexnine_unit_1954(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11232)
);

ninexnine_unit ninexnine_unit_1955(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12232)
);

assign C1232=c10232+c11232+c12232;
assign A1232=(C1232>=0)?1:0;

assign P2232=A1232;

ninexnine_unit ninexnine_unit_1956(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10242)
);

ninexnine_unit ninexnine_unit_1957(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11242)
);

ninexnine_unit ninexnine_unit_1958(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12242)
);

assign C1242=c10242+c11242+c12242;
assign A1242=(C1242>=0)?1:0;

assign P2242=A1242;

ninexnine_unit ninexnine_unit_1959(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10302)
);

ninexnine_unit ninexnine_unit_1960(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11302)
);

ninexnine_unit ninexnine_unit_1961(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12302)
);

assign C1302=c10302+c11302+c12302;
assign A1302=(C1302>=0)?1:0;

assign P2302=A1302;

ninexnine_unit ninexnine_unit_1962(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10312)
);

ninexnine_unit ninexnine_unit_1963(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11312)
);

ninexnine_unit ninexnine_unit_1964(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12312)
);

assign C1312=c10312+c11312+c12312;
assign A1312=(C1312>=0)?1:0;

assign P2312=A1312;

ninexnine_unit ninexnine_unit_1965(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10322)
);

ninexnine_unit ninexnine_unit_1966(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11322)
);

ninexnine_unit ninexnine_unit_1967(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12322)
);

assign C1322=c10322+c11322+c12322;
assign A1322=(C1322>=0)?1:0;

assign P2322=A1322;

ninexnine_unit ninexnine_unit_1968(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10332)
);

ninexnine_unit ninexnine_unit_1969(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11332)
);

ninexnine_unit ninexnine_unit_1970(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12332)
);

assign C1332=c10332+c11332+c12332;
assign A1332=(C1332>=0)?1:0;

assign P2332=A1332;

ninexnine_unit ninexnine_unit_1971(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10342)
);

ninexnine_unit ninexnine_unit_1972(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11342)
);

ninexnine_unit ninexnine_unit_1973(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12342)
);

assign C1342=c10342+c11342+c12342;
assign A1342=(C1342>=0)?1:0;

assign P2342=A1342;

ninexnine_unit ninexnine_unit_1974(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10402)
);

ninexnine_unit ninexnine_unit_1975(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11402)
);

ninexnine_unit ninexnine_unit_1976(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12402)
);

assign C1402=c10402+c11402+c12402;
assign A1402=(C1402>=0)?1:0;

assign P2402=A1402;

ninexnine_unit ninexnine_unit_1977(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10412)
);

ninexnine_unit ninexnine_unit_1978(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11412)
);

ninexnine_unit ninexnine_unit_1979(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12412)
);

assign C1412=c10412+c11412+c12412;
assign A1412=(C1412>=0)?1:0;

assign P2412=A1412;

ninexnine_unit ninexnine_unit_1980(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10422)
);

ninexnine_unit ninexnine_unit_1981(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11422)
);

ninexnine_unit ninexnine_unit_1982(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12422)
);

assign C1422=c10422+c11422+c12422;
assign A1422=(C1422>=0)?1:0;

assign P2422=A1422;

ninexnine_unit ninexnine_unit_1983(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10432)
);

ninexnine_unit ninexnine_unit_1984(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11432)
);

ninexnine_unit ninexnine_unit_1985(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12432)
);

assign C1432=c10432+c11432+c12432;
assign A1432=(C1432>=0)?1:0;

assign P2432=A1432;

ninexnine_unit ninexnine_unit_1986(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W12000),
				.b1(W12010),
				.b2(W12020),
				.b3(W12100),
				.b4(W12110),
				.b5(W12120),
				.b6(W12200),
				.b7(W12210),
				.b8(W12220),
				.c(c10442)
);

ninexnine_unit ninexnine_unit_1987(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W12001),
				.b1(W12011),
				.b2(W12021),
				.b3(W12101),
				.b4(W12111),
				.b5(W12121),
				.b6(W12201),
				.b7(W12211),
				.b8(W12221),
				.c(c11442)
);

ninexnine_unit ninexnine_unit_1988(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W12002),
				.b1(W12012),
				.b2(W12022),
				.b3(W12102),
				.b4(W12112),
				.b5(W12122),
				.b6(W12202),
				.b7(W12212),
				.b8(W12222),
				.c(c12442)
);

assign C1442=c10442+c11442+c12442;
assign A1442=(C1442>=0)?1:0;

assign P2442=A1442;

ninexnine_unit ninexnine_unit_1989(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10003)
);

ninexnine_unit ninexnine_unit_1990(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11003)
);

ninexnine_unit ninexnine_unit_1991(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12003)
);

assign C1003=c10003+c11003+c12003;
assign A1003=(C1003>=0)?1:0;

assign P2003=A1003;

ninexnine_unit ninexnine_unit_1992(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10013)
);

ninexnine_unit ninexnine_unit_1993(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11013)
);

ninexnine_unit ninexnine_unit_1994(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12013)
);

assign C1013=c10013+c11013+c12013;
assign A1013=(C1013>=0)?1:0;

assign P2013=A1013;

ninexnine_unit ninexnine_unit_1995(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10023)
);

ninexnine_unit ninexnine_unit_1996(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11023)
);

ninexnine_unit ninexnine_unit_1997(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12023)
);

assign C1023=c10023+c11023+c12023;
assign A1023=(C1023>=0)?1:0;

assign P2023=A1023;

ninexnine_unit ninexnine_unit_1998(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10033)
);

ninexnine_unit ninexnine_unit_1999(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11033)
);

ninexnine_unit ninexnine_unit_2000(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12033)
);

assign C1033=c10033+c11033+c12033;
assign A1033=(C1033>=0)?1:0;

assign P2033=A1033;

ninexnine_unit ninexnine_unit_2001(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10043)
);

ninexnine_unit ninexnine_unit_2002(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11043)
);

ninexnine_unit ninexnine_unit_2003(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12043)
);

assign C1043=c10043+c11043+c12043;
assign A1043=(C1043>=0)?1:0;

assign P2043=A1043;

ninexnine_unit ninexnine_unit_2004(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10103)
);

ninexnine_unit ninexnine_unit_2005(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11103)
);

ninexnine_unit ninexnine_unit_2006(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12103)
);

assign C1103=c10103+c11103+c12103;
assign A1103=(C1103>=0)?1:0;

assign P2103=A1103;

ninexnine_unit ninexnine_unit_2007(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10113)
);

ninexnine_unit ninexnine_unit_2008(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11113)
);

ninexnine_unit ninexnine_unit_2009(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12113)
);

assign C1113=c10113+c11113+c12113;
assign A1113=(C1113>=0)?1:0;

assign P2113=A1113;

ninexnine_unit ninexnine_unit_2010(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10123)
);

ninexnine_unit ninexnine_unit_2011(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11123)
);

ninexnine_unit ninexnine_unit_2012(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12123)
);

assign C1123=c10123+c11123+c12123;
assign A1123=(C1123>=0)?1:0;

assign P2123=A1123;

ninexnine_unit ninexnine_unit_2013(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10133)
);

ninexnine_unit ninexnine_unit_2014(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11133)
);

ninexnine_unit ninexnine_unit_2015(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12133)
);

assign C1133=c10133+c11133+c12133;
assign A1133=(C1133>=0)?1:0;

assign P2133=A1133;

ninexnine_unit ninexnine_unit_2016(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10143)
);

ninexnine_unit ninexnine_unit_2017(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11143)
);

ninexnine_unit ninexnine_unit_2018(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12143)
);

assign C1143=c10143+c11143+c12143;
assign A1143=(C1143>=0)?1:0;

assign P2143=A1143;

ninexnine_unit ninexnine_unit_2019(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10203)
);

ninexnine_unit ninexnine_unit_2020(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11203)
);

ninexnine_unit ninexnine_unit_2021(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12203)
);

assign C1203=c10203+c11203+c12203;
assign A1203=(C1203>=0)?1:0;

assign P2203=A1203;

ninexnine_unit ninexnine_unit_2022(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10213)
);

ninexnine_unit ninexnine_unit_2023(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11213)
);

ninexnine_unit ninexnine_unit_2024(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12213)
);

assign C1213=c10213+c11213+c12213;
assign A1213=(C1213>=0)?1:0;

assign P2213=A1213;

ninexnine_unit ninexnine_unit_2025(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10223)
);

ninexnine_unit ninexnine_unit_2026(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11223)
);

ninexnine_unit ninexnine_unit_2027(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12223)
);

assign C1223=c10223+c11223+c12223;
assign A1223=(C1223>=0)?1:0;

assign P2223=A1223;

ninexnine_unit ninexnine_unit_2028(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10233)
);

ninexnine_unit ninexnine_unit_2029(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11233)
);

ninexnine_unit ninexnine_unit_2030(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12233)
);

assign C1233=c10233+c11233+c12233;
assign A1233=(C1233>=0)?1:0;

assign P2233=A1233;

ninexnine_unit ninexnine_unit_2031(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10243)
);

ninexnine_unit ninexnine_unit_2032(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11243)
);

ninexnine_unit ninexnine_unit_2033(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12243)
);

assign C1243=c10243+c11243+c12243;
assign A1243=(C1243>=0)?1:0;

assign P2243=A1243;

ninexnine_unit ninexnine_unit_2034(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10303)
);

ninexnine_unit ninexnine_unit_2035(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11303)
);

ninexnine_unit ninexnine_unit_2036(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12303)
);

assign C1303=c10303+c11303+c12303;
assign A1303=(C1303>=0)?1:0;

assign P2303=A1303;

ninexnine_unit ninexnine_unit_2037(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10313)
);

ninexnine_unit ninexnine_unit_2038(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11313)
);

ninexnine_unit ninexnine_unit_2039(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12313)
);

assign C1313=c10313+c11313+c12313;
assign A1313=(C1313>=0)?1:0;

assign P2313=A1313;

ninexnine_unit ninexnine_unit_2040(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10323)
);

ninexnine_unit ninexnine_unit_2041(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11323)
);

ninexnine_unit ninexnine_unit_2042(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12323)
);

assign C1323=c10323+c11323+c12323;
assign A1323=(C1323>=0)?1:0;

assign P2323=A1323;

ninexnine_unit ninexnine_unit_2043(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10333)
);

ninexnine_unit ninexnine_unit_2044(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11333)
);

ninexnine_unit ninexnine_unit_2045(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12333)
);

assign C1333=c10333+c11333+c12333;
assign A1333=(C1333>=0)?1:0;

assign P2333=A1333;

ninexnine_unit ninexnine_unit_2046(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10343)
);

ninexnine_unit ninexnine_unit_2047(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11343)
);

ninexnine_unit ninexnine_unit_2048(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12343)
);

assign C1343=c10343+c11343+c12343;
assign A1343=(C1343>=0)?1:0;

assign P2343=A1343;

ninexnine_unit ninexnine_unit_2049(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10403)
);

ninexnine_unit ninexnine_unit_2050(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11403)
);

ninexnine_unit ninexnine_unit_2051(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12403)
);

assign C1403=c10403+c11403+c12403;
assign A1403=(C1403>=0)?1:0;

assign P2403=A1403;

ninexnine_unit ninexnine_unit_2052(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10413)
);

ninexnine_unit ninexnine_unit_2053(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11413)
);

ninexnine_unit ninexnine_unit_2054(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12413)
);

assign C1413=c10413+c11413+c12413;
assign A1413=(C1413>=0)?1:0;

assign P2413=A1413;

ninexnine_unit ninexnine_unit_2055(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10423)
);

ninexnine_unit ninexnine_unit_2056(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11423)
);

ninexnine_unit ninexnine_unit_2057(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12423)
);

assign C1423=c10423+c11423+c12423;
assign A1423=(C1423>=0)?1:0;

assign P2423=A1423;

ninexnine_unit ninexnine_unit_2058(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10433)
);

ninexnine_unit ninexnine_unit_2059(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11433)
);

ninexnine_unit ninexnine_unit_2060(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12433)
);

assign C1433=c10433+c11433+c12433;
assign A1433=(C1433>=0)?1:0;

assign P2433=A1433;

ninexnine_unit ninexnine_unit_2061(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W13000),
				.b1(W13010),
				.b2(W13020),
				.b3(W13100),
				.b4(W13110),
				.b5(W13120),
				.b6(W13200),
				.b7(W13210),
				.b8(W13220),
				.c(c10443)
);

ninexnine_unit ninexnine_unit_2062(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W13001),
				.b1(W13011),
				.b2(W13021),
				.b3(W13101),
				.b4(W13111),
				.b5(W13121),
				.b6(W13201),
				.b7(W13211),
				.b8(W13221),
				.c(c11443)
);

ninexnine_unit ninexnine_unit_2063(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W13002),
				.b1(W13012),
				.b2(W13022),
				.b3(W13102),
				.b4(W13112),
				.b5(W13122),
				.b6(W13202),
				.b7(W13212),
				.b8(W13222),
				.c(c12443)
);

assign C1443=c10443+c11443+c12443;
assign A1443=(C1443>=0)?1:0;

assign P2443=A1443;

ninexnine_unit ninexnine_unit_2064(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10004)
);

ninexnine_unit ninexnine_unit_2065(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11004)
);

ninexnine_unit ninexnine_unit_2066(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12004)
);

assign C1004=c10004+c11004+c12004;
assign A1004=(C1004>=0)?1:0;

assign P2004=A1004;

ninexnine_unit ninexnine_unit_2067(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10014)
);

ninexnine_unit ninexnine_unit_2068(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11014)
);

ninexnine_unit ninexnine_unit_2069(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12014)
);

assign C1014=c10014+c11014+c12014;
assign A1014=(C1014>=0)?1:0;

assign P2014=A1014;

ninexnine_unit ninexnine_unit_2070(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10024)
);

ninexnine_unit ninexnine_unit_2071(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11024)
);

ninexnine_unit ninexnine_unit_2072(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12024)
);

assign C1024=c10024+c11024+c12024;
assign A1024=(C1024>=0)?1:0;

assign P2024=A1024;

ninexnine_unit ninexnine_unit_2073(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10034)
);

ninexnine_unit ninexnine_unit_2074(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11034)
);

ninexnine_unit ninexnine_unit_2075(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12034)
);

assign C1034=c10034+c11034+c12034;
assign A1034=(C1034>=0)?1:0;

assign P2034=A1034;

ninexnine_unit ninexnine_unit_2076(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10044)
);

ninexnine_unit ninexnine_unit_2077(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11044)
);

ninexnine_unit ninexnine_unit_2078(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12044)
);

assign C1044=c10044+c11044+c12044;
assign A1044=(C1044>=0)?1:0;

assign P2044=A1044;

ninexnine_unit ninexnine_unit_2079(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10104)
);

ninexnine_unit ninexnine_unit_2080(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11104)
);

ninexnine_unit ninexnine_unit_2081(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12104)
);

assign C1104=c10104+c11104+c12104;
assign A1104=(C1104>=0)?1:0;

assign P2104=A1104;

ninexnine_unit ninexnine_unit_2082(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10114)
);

ninexnine_unit ninexnine_unit_2083(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11114)
);

ninexnine_unit ninexnine_unit_2084(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12114)
);

assign C1114=c10114+c11114+c12114;
assign A1114=(C1114>=0)?1:0;

assign P2114=A1114;

ninexnine_unit ninexnine_unit_2085(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10124)
);

ninexnine_unit ninexnine_unit_2086(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11124)
);

ninexnine_unit ninexnine_unit_2087(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12124)
);

assign C1124=c10124+c11124+c12124;
assign A1124=(C1124>=0)?1:0;

assign P2124=A1124;

ninexnine_unit ninexnine_unit_2088(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10134)
);

ninexnine_unit ninexnine_unit_2089(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11134)
);

ninexnine_unit ninexnine_unit_2090(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12134)
);

assign C1134=c10134+c11134+c12134;
assign A1134=(C1134>=0)?1:0;

assign P2134=A1134;

ninexnine_unit ninexnine_unit_2091(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10144)
);

ninexnine_unit ninexnine_unit_2092(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11144)
);

ninexnine_unit ninexnine_unit_2093(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12144)
);

assign C1144=c10144+c11144+c12144;
assign A1144=(C1144>=0)?1:0;

assign P2144=A1144;

ninexnine_unit ninexnine_unit_2094(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10204)
);

ninexnine_unit ninexnine_unit_2095(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11204)
);

ninexnine_unit ninexnine_unit_2096(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12204)
);

assign C1204=c10204+c11204+c12204;
assign A1204=(C1204>=0)?1:0;

assign P2204=A1204;

ninexnine_unit ninexnine_unit_2097(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10214)
);

ninexnine_unit ninexnine_unit_2098(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11214)
);

ninexnine_unit ninexnine_unit_2099(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12214)
);

assign C1214=c10214+c11214+c12214;
assign A1214=(C1214>=0)?1:0;

assign P2214=A1214;

ninexnine_unit ninexnine_unit_2100(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10224)
);

ninexnine_unit ninexnine_unit_2101(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11224)
);

ninexnine_unit ninexnine_unit_2102(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12224)
);

assign C1224=c10224+c11224+c12224;
assign A1224=(C1224>=0)?1:0;

assign P2224=A1224;

ninexnine_unit ninexnine_unit_2103(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10234)
);

ninexnine_unit ninexnine_unit_2104(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11234)
);

ninexnine_unit ninexnine_unit_2105(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12234)
);

assign C1234=c10234+c11234+c12234;
assign A1234=(C1234>=0)?1:0;

assign P2234=A1234;

ninexnine_unit ninexnine_unit_2106(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10244)
);

ninexnine_unit ninexnine_unit_2107(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11244)
);

ninexnine_unit ninexnine_unit_2108(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12244)
);

assign C1244=c10244+c11244+c12244;
assign A1244=(C1244>=0)?1:0;

assign P2244=A1244;

ninexnine_unit ninexnine_unit_2109(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10304)
);

ninexnine_unit ninexnine_unit_2110(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11304)
);

ninexnine_unit ninexnine_unit_2111(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12304)
);

assign C1304=c10304+c11304+c12304;
assign A1304=(C1304>=0)?1:0;

assign P2304=A1304;

ninexnine_unit ninexnine_unit_2112(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10314)
);

ninexnine_unit ninexnine_unit_2113(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11314)
);

ninexnine_unit ninexnine_unit_2114(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12314)
);

assign C1314=c10314+c11314+c12314;
assign A1314=(C1314>=0)?1:0;

assign P2314=A1314;

ninexnine_unit ninexnine_unit_2115(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10324)
);

ninexnine_unit ninexnine_unit_2116(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11324)
);

ninexnine_unit ninexnine_unit_2117(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12324)
);

assign C1324=c10324+c11324+c12324;
assign A1324=(C1324>=0)?1:0;

assign P2324=A1324;

ninexnine_unit ninexnine_unit_2118(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10334)
);

ninexnine_unit ninexnine_unit_2119(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11334)
);

ninexnine_unit ninexnine_unit_2120(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12334)
);

assign C1334=c10334+c11334+c12334;
assign A1334=(C1334>=0)?1:0;

assign P2334=A1334;

ninexnine_unit ninexnine_unit_2121(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10344)
);

ninexnine_unit ninexnine_unit_2122(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11344)
);

ninexnine_unit ninexnine_unit_2123(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12344)
);

assign C1344=c10344+c11344+c12344;
assign A1344=(C1344>=0)?1:0;

assign P2344=A1344;

ninexnine_unit ninexnine_unit_2124(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10404)
);

ninexnine_unit ninexnine_unit_2125(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11404)
);

ninexnine_unit ninexnine_unit_2126(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12404)
);

assign C1404=c10404+c11404+c12404;
assign A1404=(C1404>=0)?1:0;

assign P2404=A1404;

ninexnine_unit ninexnine_unit_2127(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10414)
);

ninexnine_unit ninexnine_unit_2128(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11414)
);

ninexnine_unit ninexnine_unit_2129(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12414)
);

assign C1414=c10414+c11414+c12414;
assign A1414=(C1414>=0)?1:0;

assign P2414=A1414;

ninexnine_unit ninexnine_unit_2130(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10424)
);

ninexnine_unit ninexnine_unit_2131(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11424)
);

ninexnine_unit ninexnine_unit_2132(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12424)
);

assign C1424=c10424+c11424+c12424;
assign A1424=(C1424>=0)?1:0;

assign P2424=A1424;

ninexnine_unit ninexnine_unit_2133(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10434)
);

ninexnine_unit ninexnine_unit_2134(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11434)
);

ninexnine_unit ninexnine_unit_2135(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12434)
);

assign C1434=c10434+c11434+c12434;
assign A1434=(C1434>=0)?1:0;

assign P2434=A1434;

ninexnine_unit ninexnine_unit_2136(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W14000),
				.b1(W14010),
				.b2(W14020),
				.b3(W14100),
				.b4(W14110),
				.b5(W14120),
				.b6(W14200),
				.b7(W14210),
				.b8(W14220),
				.c(c10444)
);

ninexnine_unit ninexnine_unit_2137(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W14001),
				.b1(W14011),
				.b2(W14021),
				.b3(W14101),
				.b4(W14111),
				.b5(W14121),
				.b6(W14201),
				.b7(W14211),
				.b8(W14221),
				.c(c11444)
);

ninexnine_unit ninexnine_unit_2138(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W14002),
				.b1(W14012),
				.b2(W14022),
				.b3(W14102),
				.b4(W14112),
				.b5(W14122),
				.b6(W14202),
				.b7(W14212),
				.b8(W14222),
				.c(c12444)
);

assign C1444=c10444+c11444+c12444;
assign A1444=(C1444>=0)?1:0;

assign P2444=A1444;

ninexnine_unit ninexnine_unit_2139(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10005)
);

ninexnine_unit ninexnine_unit_2140(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11005)
);

ninexnine_unit ninexnine_unit_2141(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12005)
);

assign C1005=c10005+c11005+c12005;
assign A1005=(C1005>=0)?1:0;

assign P2005=A1005;

ninexnine_unit ninexnine_unit_2142(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10015)
);

ninexnine_unit ninexnine_unit_2143(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11015)
);

ninexnine_unit ninexnine_unit_2144(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12015)
);

assign C1015=c10015+c11015+c12015;
assign A1015=(C1015>=0)?1:0;

assign P2015=A1015;

ninexnine_unit ninexnine_unit_2145(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10025)
);

ninexnine_unit ninexnine_unit_2146(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11025)
);

ninexnine_unit ninexnine_unit_2147(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12025)
);

assign C1025=c10025+c11025+c12025;
assign A1025=(C1025>=0)?1:0;

assign P2025=A1025;

ninexnine_unit ninexnine_unit_2148(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10035)
);

ninexnine_unit ninexnine_unit_2149(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11035)
);

ninexnine_unit ninexnine_unit_2150(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12035)
);

assign C1035=c10035+c11035+c12035;
assign A1035=(C1035>=0)?1:0;

assign P2035=A1035;

ninexnine_unit ninexnine_unit_2151(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10045)
);

ninexnine_unit ninexnine_unit_2152(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11045)
);

ninexnine_unit ninexnine_unit_2153(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12045)
);

assign C1045=c10045+c11045+c12045;
assign A1045=(C1045>=0)?1:0;

assign P2045=A1045;

ninexnine_unit ninexnine_unit_2154(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10105)
);

ninexnine_unit ninexnine_unit_2155(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11105)
);

ninexnine_unit ninexnine_unit_2156(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12105)
);

assign C1105=c10105+c11105+c12105;
assign A1105=(C1105>=0)?1:0;

assign P2105=A1105;

ninexnine_unit ninexnine_unit_2157(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10115)
);

ninexnine_unit ninexnine_unit_2158(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11115)
);

ninexnine_unit ninexnine_unit_2159(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12115)
);

assign C1115=c10115+c11115+c12115;
assign A1115=(C1115>=0)?1:0;

assign P2115=A1115;

ninexnine_unit ninexnine_unit_2160(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10125)
);

ninexnine_unit ninexnine_unit_2161(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11125)
);

ninexnine_unit ninexnine_unit_2162(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12125)
);

assign C1125=c10125+c11125+c12125;
assign A1125=(C1125>=0)?1:0;

assign P2125=A1125;

ninexnine_unit ninexnine_unit_2163(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10135)
);

ninexnine_unit ninexnine_unit_2164(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11135)
);

ninexnine_unit ninexnine_unit_2165(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12135)
);

assign C1135=c10135+c11135+c12135;
assign A1135=(C1135>=0)?1:0;

assign P2135=A1135;

ninexnine_unit ninexnine_unit_2166(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10145)
);

ninexnine_unit ninexnine_unit_2167(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11145)
);

ninexnine_unit ninexnine_unit_2168(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12145)
);

assign C1145=c10145+c11145+c12145;
assign A1145=(C1145>=0)?1:0;

assign P2145=A1145;

ninexnine_unit ninexnine_unit_2169(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10205)
);

ninexnine_unit ninexnine_unit_2170(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11205)
);

ninexnine_unit ninexnine_unit_2171(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12205)
);

assign C1205=c10205+c11205+c12205;
assign A1205=(C1205>=0)?1:0;

assign P2205=A1205;

ninexnine_unit ninexnine_unit_2172(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10215)
);

ninexnine_unit ninexnine_unit_2173(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11215)
);

ninexnine_unit ninexnine_unit_2174(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12215)
);

assign C1215=c10215+c11215+c12215;
assign A1215=(C1215>=0)?1:0;

assign P2215=A1215;

ninexnine_unit ninexnine_unit_2175(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10225)
);

ninexnine_unit ninexnine_unit_2176(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11225)
);

ninexnine_unit ninexnine_unit_2177(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12225)
);

assign C1225=c10225+c11225+c12225;
assign A1225=(C1225>=0)?1:0;

assign P2225=A1225;

ninexnine_unit ninexnine_unit_2178(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10235)
);

ninexnine_unit ninexnine_unit_2179(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11235)
);

ninexnine_unit ninexnine_unit_2180(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12235)
);

assign C1235=c10235+c11235+c12235;
assign A1235=(C1235>=0)?1:0;

assign P2235=A1235;

ninexnine_unit ninexnine_unit_2181(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10245)
);

ninexnine_unit ninexnine_unit_2182(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11245)
);

ninexnine_unit ninexnine_unit_2183(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12245)
);

assign C1245=c10245+c11245+c12245;
assign A1245=(C1245>=0)?1:0;

assign P2245=A1245;

ninexnine_unit ninexnine_unit_2184(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10305)
);

ninexnine_unit ninexnine_unit_2185(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11305)
);

ninexnine_unit ninexnine_unit_2186(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12305)
);

assign C1305=c10305+c11305+c12305;
assign A1305=(C1305>=0)?1:0;

assign P2305=A1305;

ninexnine_unit ninexnine_unit_2187(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10315)
);

ninexnine_unit ninexnine_unit_2188(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11315)
);

ninexnine_unit ninexnine_unit_2189(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12315)
);

assign C1315=c10315+c11315+c12315;
assign A1315=(C1315>=0)?1:0;

assign P2315=A1315;

ninexnine_unit ninexnine_unit_2190(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10325)
);

ninexnine_unit ninexnine_unit_2191(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11325)
);

ninexnine_unit ninexnine_unit_2192(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12325)
);

assign C1325=c10325+c11325+c12325;
assign A1325=(C1325>=0)?1:0;

assign P2325=A1325;

ninexnine_unit ninexnine_unit_2193(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10335)
);

ninexnine_unit ninexnine_unit_2194(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11335)
);

ninexnine_unit ninexnine_unit_2195(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12335)
);

assign C1335=c10335+c11335+c12335;
assign A1335=(C1335>=0)?1:0;

assign P2335=A1335;

ninexnine_unit ninexnine_unit_2196(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10345)
);

ninexnine_unit ninexnine_unit_2197(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11345)
);

ninexnine_unit ninexnine_unit_2198(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12345)
);

assign C1345=c10345+c11345+c12345;
assign A1345=(C1345>=0)?1:0;

assign P2345=A1345;

ninexnine_unit ninexnine_unit_2199(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10405)
);

ninexnine_unit ninexnine_unit_2200(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11405)
);

ninexnine_unit ninexnine_unit_2201(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12405)
);

assign C1405=c10405+c11405+c12405;
assign A1405=(C1405>=0)?1:0;

assign P2405=A1405;

ninexnine_unit ninexnine_unit_2202(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10415)
);

ninexnine_unit ninexnine_unit_2203(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11415)
);

ninexnine_unit ninexnine_unit_2204(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12415)
);

assign C1415=c10415+c11415+c12415;
assign A1415=(C1415>=0)?1:0;

assign P2415=A1415;

ninexnine_unit ninexnine_unit_2205(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10425)
);

ninexnine_unit ninexnine_unit_2206(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11425)
);

ninexnine_unit ninexnine_unit_2207(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12425)
);

assign C1425=c10425+c11425+c12425;
assign A1425=(C1425>=0)?1:0;

assign P2425=A1425;

ninexnine_unit ninexnine_unit_2208(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10435)
);

ninexnine_unit ninexnine_unit_2209(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11435)
);

ninexnine_unit ninexnine_unit_2210(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12435)
);

assign C1435=c10435+c11435+c12435;
assign A1435=(C1435>=0)?1:0;

assign P2435=A1435;

ninexnine_unit ninexnine_unit_2211(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W15000),
				.b1(W15010),
				.b2(W15020),
				.b3(W15100),
				.b4(W15110),
				.b5(W15120),
				.b6(W15200),
				.b7(W15210),
				.b8(W15220),
				.c(c10445)
);

ninexnine_unit ninexnine_unit_2212(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W15001),
				.b1(W15011),
				.b2(W15021),
				.b3(W15101),
				.b4(W15111),
				.b5(W15121),
				.b6(W15201),
				.b7(W15211),
				.b8(W15221),
				.c(c11445)
);

ninexnine_unit ninexnine_unit_2213(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W15002),
				.b1(W15012),
				.b2(W15022),
				.b3(W15102),
				.b4(W15112),
				.b5(W15122),
				.b6(W15202),
				.b7(W15212),
				.b8(W15222),
				.c(c12445)
);

assign C1445=c10445+c11445+c12445;
assign A1445=(C1445>=0)?1:0;

assign P2445=A1445;

ninexnine_unit ninexnine_unit_2214(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10006)
);

ninexnine_unit ninexnine_unit_2215(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11006)
);

ninexnine_unit ninexnine_unit_2216(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12006)
);

assign C1006=c10006+c11006+c12006;
assign A1006=(C1006>=0)?1:0;

assign P2006=A1006;

ninexnine_unit ninexnine_unit_2217(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10016)
);

ninexnine_unit ninexnine_unit_2218(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11016)
);

ninexnine_unit ninexnine_unit_2219(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12016)
);

assign C1016=c10016+c11016+c12016;
assign A1016=(C1016>=0)?1:0;

assign P2016=A1016;

ninexnine_unit ninexnine_unit_2220(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10026)
);

ninexnine_unit ninexnine_unit_2221(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11026)
);

ninexnine_unit ninexnine_unit_2222(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12026)
);

assign C1026=c10026+c11026+c12026;
assign A1026=(C1026>=0)?1:0;

assign P2026=A1026;

ninexnine_unit ninexnine_unit_2223(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10036)
);

ninexnine_unit ninexnine_unit_2224(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11036)
);

ninexnine_unit ninexnine_unit_2225(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12036)
);

assign C1036=c10036+c11036+c12036;
assign A1036=(C1036>=0)?1:0;

assign P2036=A1036;

ninexnine_unit ninexnine_unit_2226(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10046)
);

ninexnine_unit ninexnine_unit_2227(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11046)
);

ninexnine_unit ninexnine_unit_2228(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12046)
);

assign C1046=c10046+c11046+c12046;
assign A1046=(C1046>=0)?1:0;

assign P2046=A1046;

ninexnine_unit ninexnine_unit_2229(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10106)
);

ninexnine_unit ninexnine_unit_2230(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11106)
);

ninexnine_unit ninexnine_unit_2231(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12106)
);

assign C1106=c10106+c11106+c12106;
assign A1106=(C1106>=0)?1:0;

assign P2106=A1106;

ninexnine_unit ninexnine_unit_2232(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10116)
);

ninexnine_unit ninexnine_unit_2233(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11116)
);

ninexnine_unit ninexnine_unit_2234(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12116)
);

assign C1116=c10116+c11116+c12116;
assign A1116=(C1116>=0)?1:0;

assign P2116=A1116;

ninexnine_unit ninexnine_unit_2235(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10126)
);

ninexnine_unit ninexnine_unit_2236(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11126)
);

ninexnine_unit ninexnine_unit_2237(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12126)
);

assign C1126=c10126+c11126+c12126;
assign A1126=(C1126>=0)?1:0;

assign P2126=A1126;

ninexnine_unit ninexnine_unit_2238(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10136)
);

ninexnine_unit ninexnine_unit_2239(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11136)
);

ninexnine_unit ninexnine_unit_2240(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12136)
);

assign C1136=c10136+c11136+c12136;
assign A1136=(C1136>=0)?1:0;

assign P2136=A1136;

ninexnine_unit ninexnine_unit_2241(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10146)
);

ninexnine_unit ninexnine_unit_2242(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11146)
);

ninexnine_unit ninexnine_unit_2243(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12146)
);

assign C1146=c10146+c11146+c12146;
assign A1146=(C1146>=0)?1:0;

assign P2146=A1146;

ninexnine_unit ninexnine_unit_2244(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10206)
);

ninexnine_unit ninexnine_unit_2245(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11206)
);

ninexnine_unit ninexnine_unit_2246(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12206)
);

assign C1206=c10206+c11206+c12206;
assign A1206=(C1206>=0)?1:0;

assign P2206=A1206;

ninexnine_unit ninexnine_unit_2247(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10216)
);

ninexnine_unit ninexnine_unit_2248(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11216)
);

ninexnine_unit ninexnine_unit_2249(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12216)
);

assign C1216=c10216+c11216+c12216;
assign A1216=(C1216>=0)?1:0;

assign P2216=A1216;

ninexnine_unit ninexnine_unit_2250(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10226)
);

ninexnine_unit ninexnine_unit_2251(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11226)
);

ninexnine_unit ninexnine_unit_2252(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12226)
);

assign C1226=c10226+c11226+c12226;
assign A1226=(C1226>=0)?1:0;

assign P2226=A1226;

ninexnine_unit ninexnine_unit_2253(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10236)
);

ninexnine_unit ninexnine_unit_2254(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11236)
);

ninexnine_unit ninexnine_unit_2255(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12236)
);

assign C1236=c10236+c11236+c12236;
assign A1236=(C1236>=0)?1:0;

assign P2236=A1236;

ninexnine_unit ninexnine_unit_2256(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10246)
);

ninexnine_unit ninexnine_unit_2257(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11246)
);

ninexnine_unit ninexnine_unit_2258(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12246)
);

assign C1246=c10246+c11246+c12246;
assign A1246=(C1246>=0)?1:0;

assign P2246=A1246;

ninexnine_unit ninexnine_unit_2259(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10306)
);

ninexnine_unit ninexnine_unit_2260(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11306)
);

ninexnine_unit ninexnine_unit_2261(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12306)
);

assign C1306=c10306+c11306+c12306;
assign A1306=(C1306>=0)?1:0;

assign P2306=A1306;

ninexnine_unit ninexnine_unit_2262(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10316)
);

ninexnine_unit ninexnine_unit_2263(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11316)
);

ninexnine_unit ninexnine_unit_2264(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12316)
);

assign C1316=c10316+c11316+c12316;
assign A1316=(C1316>=0)?1:0;

assign P2316=A1316;

ninexnine_unit ninexnine_unit_2265(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10326)
);

ninexnine_unit ninexnine_unit_2266(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11326)
);

ninexnine_unit ninexnine_unit_2267(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12326)
);

assign C1326=c10326+c11326+c12326;
assign A1326=(C1326>=0)?1:0;

assign P2326=A1326;

ninexnine_unit ninexnine_unit_2268(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10336)
);

ninexnine_unit ninexnine_unit_2269(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11336)
);

ninexnine_unit ninexnine_unit_2270(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12336)
);

assign C1336=c10336+c11336+c12336;
assign A1336=(C1336>=0)?1:0;

assign P2336=A1336;

ninexnine_unit ninexnine_unit_2271(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10346)
);

ninexnine_unit ninexnine_unit_2272(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11346)
);

ninexnine_unit ninexnine_unit_2273(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12346)
);

assign C1346=c10346+c11346+c12346;
assign A1346=(C1346>=0)?1:0;

assign P2346=A1346;

ninexnine_unit ninexnine_unit_2274(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10406)
);

ninexnine_unit ninexnine_unit_2275(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11406)
);

ninexnine_unit ninexnine_unit_2276(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12406)
);

assign C1406=c10406+c11406+c12406;
assign A1406=(C1406>=0)?1:0;

assign P2406=A1406;

ninexnine_unit ninexnine_unit_2277(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10416)
);

ninexnine_unit ninexnine_unit_2278(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11416)
);

ninexnine_unit ninexnine_unit_2279(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12416)
);

assign C1416=c10416+c11416+c12416;
assign A1416=(C1416>=0)?1:0;

assign P2416=A1416;

ninexnine_unit ninexnine_unit_2280(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10426)
);

ninexnine_unit ninexnine_unit_2281(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11426)
);

ninexnine_unit ninexnine_unit_2282(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12426)
);

assign C1426=c10426+c11426+c12426;
assign A1426=(C1426>=0)?1:0;

assign P2426=A1426;

ninexnine_unit ninexnine_unit_2283(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10436)
);

ninexnine_unit ninexnine_unit_2284(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11436)
);

ninexnine_unit ninexnine_unit_2285(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12436)
);

assign C1436=c10436+c11436+c12436;
assign A1436=(C1436>=0)?1:0;

assign P2436=A1436;

ninexnine_unit ninexnine_unit_2286(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W16000),
				.b1(W16010),
				.b2(W16020),
				.b3(W16100),
				.b4(W16110),
				.b5(W16120),
				.b6(W16200),
				.b7(W16210),
				.b8(W16220),
				.c(c10446)
);

ninexnine_unit ninexnine_unit_2287(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W16001),
				.b1(W16011),
				.b2(W16021),
				.b3(W16101),
				.b4(W16111),
				.b5(W16121),
				.b6(W16201),
				.b7(W16211),
				.b8(W16221),
				.c(c11446)
);

ninexnine_unit ninexnine_unit_2288(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W16002),
				.b1(W16012),
				.b2(W16022),
				.b3(W16102),
				.b4(W16112),
				.b5(W16122),
				.b6(W16202),
				.b7(W16212),
				.b8(W16222),
				.c(c12446)
);

assign C1446=c10446+c11446+c12446;
assign A1446=(C1446>=0)?1:0;

assign P2446=A1446;

ninexnine_unit ninexnine_unit_2289(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10007)
);

ninexnine_unit ninexnine_unit_2290(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11007)
);

ninexnine_unit ninexnine_unit_2291(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12007)
);

assign C1007=c10007+c11007+c12007;
assign A1007=(C1007>=0)?1:0;

assign P2007=A1007;

ninexnine_unit ninexnine_unit_2292(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10017)
);

ninexnine_unit ninexnine_unit_2293(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11017)
);

ninexnine_unit ninexnine_unit_2294(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12017)
);

assign C1017=c10017+c11017+c12017;
assign A1017=(C1017>=0)?1:0;

assign P2017=A1017;

ninexnine_unit ninexnine_unit_2295(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10027)
);

ninexnine_unit ninexnine_unit_2296(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11027)
);

ninexnine_unit ninexnine_unit_2297(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12027)
);

assign C1027=c10027+c11027+c12027;
assign A1027=(C1027>=0)?1:0;

assign P2027=A1027;

ninexnine_unit ninexnine_unit_2298(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10037)
);

ninexnine_unit ninexnine_unit_2299(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11037)
);

ninexnine_unit ninexnine_unit_2300(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12037)
);

assign C1037=c10037+c11037+c12037;
assign A1037=(C1037>=0)?1:0;

assign P2037=A1037;

ninexnine_unit ninexnine_unit_2301(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10047)
);

ninexnine_unit ninexnine_unit_2302(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11047)
);

ninexnine_unit ninexnine_unit_2303(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12047)
);

assign C1047=c10047+c11047+c12047;
assign A1047=(C1047>=0)?1:0;

assign P2047=A1047;

ninexnine_unit ninexnine_unit_2304(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10107)
);

ninexnine_unit ninexnine_unit_2305(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11107)
);

ninexnine_unit ninexnine_unit_2306(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12107)
);

assign C1107=c10107+c11107+c12107;
assign A1107=(C1107>=0)?1:0;

assign P2107=A1107;

ninexnine_unit ninexnine_unit_2307(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10117)
);

ninexnine_unit ninexnine_unit_2308(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11117)
);

ninexnine_unit ninexnine_unit_2309(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12117)
);

assign C1117=c10117+c11117+c12117;
assign A1117=(C1117>=0)?1:0;

assign P2117=A1117;

ninexnine_unit ninexnine_unit_2310(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10127)
);

ninexnine_unit ninexnine_unit_2311(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11127)
);

ninexnine_unit ninexnine_unit_2312(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12127)
);

assign C1127=c10127+c11127+c12127;
assign A1127=(C1127>=0)?1:0;

assign P2127=A1127;

ninexnine_unit ninexnine_unit_2313(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10137)
);

ninexnine_unit ninexnine_unit_2314(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11137)
);

ninexnine_unit ninexnine_unit_2315(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12137)
);

assign C1137=c10137+c11137+c12137;
assign A1137=(C1137>=0)?1:0;

assign P2137=A1137;

ninexnine_unit ninexnine_unit_2316(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10147)
);

ninexnine_unit ninexnine_unit_2317(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11147)
);

ninexnine_unit ninexnine_unit_2318(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12147)
);

assign C1147=c10147+c11147+c12147;
assign A1147=(C1147>=0)?1:0;

assign P2147=A1147;

ninexnine_unit ninexnine_unit_2319(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10207)
);

ninexnine_unit ninexnine_unit_2320(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11207)
);

ninexnine_unit ninexnine_unit_2321(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12207)
);

assign C1207=c10207+c11207+c12207;
assign A1207=(C1207>=0)?1:0;

assign P2207=A1207;

ninexnine_unit ninexnine_unit_2322(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10217)
);

ninexnine_unit ninexnine_unit_2323(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11217)
);

ninexnine_unit ninexnine_unit_2324(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12217)
);

assign C1217=c10217+c11217+c12217;
assign A1217=(C1217>=0)?1:0;

assign P2217=A1217;

ninexnine_unit ninexnine_unit_2325(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10227)
);

ninexnine_unit ninexnine_unit_2326(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11227)
);

ninexnine_unit ninexnine_unit_2327(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12227)
);

assign C1227=c10227+c11227+c12227;
assign A1227=(C1227>=0)?1:0;

assign P2227=A1227;

ninexnine_unit ninexnine_unit_2328(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10237)
);

ninexnine_unit ninexnine_unit_2329(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11237)
);

ninexnine_unit ninexnine_unit_2330(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12237)
);

assign C1237=c10237+c11237+c12237;
assign A1237=(C1237>=0)?1:0;

assign P2237=A1237;

ninexnine_unit ninexnine_unit_2331(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10247)
);

ninexnine_unit ninexnine_unit_2332(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11247)
);

ninexnine_unit ninexnine_unit_2333(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12247)
);

assign C1247=c10247+c11247+c12247;
assign A1247=(C1247>=0)?1:0;

assign P2247=A1247;

ninexnine_unit ninexnine_unit_2334(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10307)
);

ninexnine_unit ninexnine_unit_2335(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11307)
);

ninexnine_unit ninexnine_unit_2336(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12307)
);

assign C1307=c10307+c11307+c12307;
assign A1307=(C1307>=0)?1:0;

assign P2307=A1307;

ninexnine_unit ninexnine_unit_2337(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10317)
);

ninexnine_unit ninexnine_unit_2338(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11317)
);

ninexnine_unit ninexnine_unit_2339(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12317)
);

assign C1317=c10317+c11317+c12317;
assign A1317=(C1317>=0)?1:0;

assign P2317=A1317;

ninexnine_unit ninexnine_unit_2340(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10327)
);

ninexnine_unit ninexnine_unit_2341(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11327)
);

ninexnine_unit ninexnine_unit_2342(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12327)
);

assign C1327=c10327+c11327+c12327;
assign A1327=(C1327>=0)?1:0;

assign P2327=A1327;

ninexnine_unit ninexnine_unit_2343(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10337)
);

ninexnine_unit ninexnine_unit_2344(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11337)
);

ninexnine_unit ninexnine_unit_2345(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12337)
);

assign C1337=c10337+c11337+c12337;
assign A1337=(C1337>=0)?1:0;

assign P2337=A1337;

ninexnine_unit ninexnine_unit_2346(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10347)
);

ninexnine_unit ninexnine_unit_2347(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11347)
);

ninexnine_unit ninexnine_unit_2348(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12347)
);

assign C1347=c10347+c11347+c12347;
assign A1347=(C1347>=0)?1:0;

assign P2347=A1347;

ninexnine_unit ninexnine_unit_2349(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10407)
);

ninexnine_unit ninexnine_unit_2350(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11407)
);

ninexnine_unit ninexnine_unit_2351(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12407)
);

assign C1407=c10407+c11407+c12407;
assign A1407=(C1407>=0)?1:0;

assign P2407=A1407;

ninexnine_unit ninexnine_unit_2352(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10417)
);

ninexnine_unit ninexnine_unit_2353(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11417)
);

ninexnine_unit ninexnine_unit_2354(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12417)
);

assign C1417=c10417+c11417+c12417;
assign A1417=(C1417>=0)?1:0;

assign P2417=A1417;

ninexnine_unit ninexnine_unit_2355(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10427)
);

ninexnine_unit ninexnine_unit_2356(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11427)
);

ninexnine_unit ninexnine_unit_2357(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12427)
);

assign C1427=c10427+c11427+c12427;
assign A1427=(C1427>=0)?1:0;

assign P2427=A1427;

ninexnine_unit ninexnine_unit_2358(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10437)
);

ninexnine_unit ninexnine_unit_2359(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11437)
);

ninexnine_unit ninexnine_unit_2360(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12437)
);

assign C1437=c10437+c11437+c12437;
assign A1437=(C1437>=0)?1:0;

assign P2437=A1437;

ninexnine_unit ninexnine_unit_2361(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W17000),
				.b1(W17010),
				.b2(W17020),
				.b3(W17100),
				.b4(W17110),
				.b5(W17120),
				.b6(W17200),
				.b7(W17210),
				.b8(W17220),
				.c(c10447)
);

ninexnine_unit ninexnine_unit_2362(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W17001),
				.b1(W17011),
				.b2(W17021),
				.b3(W17101),
				.b4(W17111),
				.b5(W17121),
				.b6(W17201),
				.b7(W17211),
				.b8(W17221),
				.c(c11447)
);

ninexnine_unit ninexnine_unit_2363(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W17002),
				.b1(W17012),
				.b2(W17022),
				.b3(W17102),
				.b4(W17112),
				.b5(W17122),
				.b6(W17202),
				.b7(W17212),
				.b8(W17222),
				.c(c12447)
);

assign C1447=c10447+c11447+c12447;
assign A1447=(C1447>=0)?1:0;

assign P2447=A1447;

ninexnine_unit ninexnine_unit_2364(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10008)
);

ninexnine_unit ninexnine_unit_2365(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11008)
);

ninexnine_unit ninexnine_unit_2366(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12008)
);

assign C1008=c10008+c11008+c12008;
assign A1008=(C1008>=0)?1:0;

assign P2008=A1008;

ninexnine_unit ninexnine_unit_2367(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10018)
);

ninexnine_unit ninexnine_unit_2368(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11018)
);

ninexnine_unit ninexnine_unit_2369(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12018)
);

assign C1018=c10018+c11018+c12018;
assign A1018=(C1018>=0)?1:0;

assign P2018=A1018;

ninexnine_unit ninexnine_unit_2370(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10028)
);

ninexnine_unit ninexnine_unit_2371(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11028)
);

ninexnine_unit ninexnine_unit_2372(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12028)
);

assign C1028=c10028+c11028+c12028;
assign A1028=(C1028>=0)?1:0;

assign P2028=A1028;

ninexnine_unit ninexnine_unit_2373(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10038)
);

ninexnine_unit ninexnine_unit_2374(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11038)
);

ninexnine_unit ninexnine_unit_2375(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12038)
);

assign C1038=c10038+c11038+c12038;
assign A1038=(C1038>=0)?1:0;

assign P2038=A1038;

ninexnine_unit ninexnine_unit_2376(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10048)
);

ninexnine_unit ninexnine_unit_2377(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11048)
);

ninexnine_unit ninexnine_unit_2378(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12048)
);

assign C1048=c10048+c11048+c12048;
assign A1048=(C1048>=0)?1:0;

assign P2048=A1048;

ninexnine_unit ninexnine_unit_2379(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10108)
);

ninexnine_unit ninexnine_unit_2380(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11108)
);

ninexnine_unit ninexnine_unit_2381(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12108)
);

assign C1108=c10108+c11108+c12108;
assign A1108=(C1108>=0)?1:0;

assign P2108=A1108;

ninexnine_unit ninexnine_unit_2382(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10118)
);

ninexnine_unit ninexnine_unit_2383(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11118)
);

ninexnine_unit ninexnine_unit_2384(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12118)
);

assign C1118=c10118+c11118+c12118;
assign A1118=(C1118>=0)?1:0;

assign P2118=A1118;

ninexnine_unit ninexnine_unit_2385(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10128)
);

ninexnine_unit ninexnine_unit_2386(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11128)
);

ninexnine_unit ninexnine_unit_2387(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12128)
);

assign C1128=c10128+c11128+c12128;
assign A1128=(C1128>=0)?1:0;

assign P2128=A1128;

ninexnine_unit ninexnine_unit_2388(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10138)
);

ninexnine_unit ninexnine_unit_2389(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11138)
);

ninexnine_unit ninexnine_unit_2390(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12138)
);

assign C1138=c10138+c11138+c12138;
assign A1138=(C1138>=0)?1:0;

assign P2138=A1138;

ninexnine_unit ninexnine_unit_2391(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10148)
);

ninexnine_unit ninexnine_unit_2392(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11148)
);

ninexnine_unit ninexnine_unit_2393(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12148)
);

assign C1148=c10148+c11148+c12148;
assign A1148=(C1148>=0)?1:0;

assign P2148=A1148;

ninexnine_unit ninexnine_unit_2394(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10208)
);

ninexnine_unit ninexnine_unit_2395(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11208)
);

ninexnine_unit ninexnine_unit_2396(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12208)
);

assign C1208=c10208+c11208+c12208;
assign A1208=(C1208>=0)?1:0;

assign P2208=A1208;

ninexnine_unit ninexnine_unit_2397(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10218)
);

ninexnine_unit ninexnine_unit_2398(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11218)
);

ninexnine_unit ninexnine_unit_2399(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12218)
);

assign C1218=c10218+c11218+c12218;
assign A1218=(C1218>=0)?1:0;

assign P2218=A1218;

ninexnine_unit ninexnine_unit_2400(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10228)
);

ninexnine_unit ninexnine_unit_2401(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11228)
);

ninexnine_unit ninexnine_unit_2402(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12228)
);

assign C1228=c10228+c11228+c12228;
assign A1228=(C1228>=0)?1:0;

assign P2228=A1228;

ninexnine_unit ninexnine_unit_2403(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10238)
);

ninexnine_unit ninexnine_unit_2404(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11238)
);

ninexnine_unit ninexnine_unit_2405(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12238)
);

assign C1238=c10238+c11238+c12238;
assign A1238=(C1238>=0)?1:0;

assign P2238=A1238;

ninexnine_unit ninexnine_unit_2406(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10248)
);

ninexnine_unit ninexnine_unit_2407(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11248)
);

ninexnine_unit ninexnine_unit_2408(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12248)
);

assign C1248=c10248+c11248+c12248;
assign A1248=(C1248>=0)?1:0;

assign P2248=A1248;

ninexnine_unit ninexnine_unit_2409(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10308)
);

ninexnine_unit ninexnine_unit_2410(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11308)
);

ninexnine_unit ninexnine_unit_2411(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12308)
);

assign C1308=c10308+c11308+c12308;
assign A1308=(C1308>=0)?1:0;

assign P2308=A1308;

ninexnine_unit ninexnine_unit_2412(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10318)
);

ninexnine_unit ninexnine_unit_2413(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11318)
);

ninexnine_unit ninexnine_unit_2414(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12318)
);

assign C1318=c10318+c11318+c12318;
assign A1318=(C1318>=0)?1:0;

assign P2318=A1318;

ninexnine_unit ninexnine_unit_2415(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10328)
);

ninexnine_unit ninexnine_unit_2416(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11328)
);

ninexnine_unit ninexnine_unit_2417(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12328)
);

assign C1328=c10328+c11328+c12328;
assign A1328=(C1328>=0)?1:0;

assign P2328=A1328;

ninexnine_unit ninexnine_unit_2418(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10338)
);

ninexnine_unit ninexnine_unit_2419(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11338)
);

ninexnine_unit ninexnine_unit_2420(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12338)
);

assign C1338=c10338+c11338+c12338;
assign A1338=(C1338>=0)?1:0;

assign P2338=A1338;

ninexnine_unit ninexnine_unit_2421(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10348)
);

ninexnine_unit ninexnine_unit_2422(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11348)
);

ninexnine_unit ninexnine_unit_2423(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12348)
);

assign C1348=c10348+c11348+c12348;
assign A1348=(C1348>=0)?1:0;

assign P2348=A1348;

ninexnine_unit ninexnine_unit_2424(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10408)
);

ninexnine_unit ninexnine_unit_2425(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11408)
);

ninexnine_unit ninexnine_unit_2426(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12408)
);

assign C1408=c10408+c11408+c12408;
assign A1408=(C1408>=0)?1:0;

assign P2408=A1408;

ninexnine_unit ninexnine_unit_2427(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10418)
);

ninexnine_unit ninexnine_unit_2428(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11418)
);

ninexnine_unit ninexnine_unit_2429(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12418)
);

assign C1418=c10418+c11418+c12418;
assign A1418=(C1418>=0)?1:0;

assign P2418=A1418;

ninexnine_unit ninexnine_unit_2430(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10428)
);

ninexnine_unit ninexnine_unit_2431(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11428)
);

ninexnine_unit ninexnine_unit_2432(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12428)
);

assign C1428=c10428+c11428+c12428;
assign A1428=(C1428>=0)?1:0;

assign P2428=A1428;

ninexnine_unit ninexnine_unit_2433(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10438)
);

ninexnine_unit ninexnine_unit_2434(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11438)
);

ninexnine_unit ninexnine_unit_2435(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12438)
);

assign C1438=c10438+c11438+c12438;
assign A1438=(C1438>=0)?1:0;

assign P2438=A1438;

ninexnine_unit ninexnine_unit_2436(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W18000),
				.b1(W18010),
				.b2(W18020),
				.b3(W18100),
				.b4(W18110),
				.b5(W18120),
				.b6(W18200),
				.b7(W18210),
				.b8(W18220),
				.c(c10448)
);

ninexnine_unit ninexnine_unit_2437(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W18001),
				.b1(W18011),
				.b2(W18021),
				.b3(W18101),
				.b4(W18111),
				.b5(W18121),
				.b6(W18201),
				.b7(W18211),
				.b8(W18221),
				.c(c11448)
);

ninexnine_unit ninexnine_unit_2438(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W18002),
				.b1(W18012),
				.b2(W18022),
				.b3(W18102),
				.b4(W18112),
				.b5(W18122),
				.b6(W18202),
				.b7(W18212),
				.b8(W18222),
				.c(c12448)
);

assign C1448=c10448+c11448+c12448;
assign A1448=(C1448>=0)?1:0;

assign P2448=A1448;

ninexnine_unit ninexnine_unit_2439(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10009)
);

ninexnine_unit ninexnine_unit_2440(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11009)
);

ninexnine_unit ninexnine_unit_2441(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12009)
);

assign C1009=c10009+c11009+c12009;
assign A1009=(C1009>=0)?1:0;

assign P2009=A1009;

ninexnine_unit ninexnine_unit_2442(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10019)
);

ninexnine_unit ninexnine_unit_2443(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11019)
);

ninexnine_unit ninexnine_unit_2444(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12019)
);

assign C1019=c10019+c11019+c12019;
assign A1019=(C1019>=0)?1:0;

assign P2019=A1019;

ninexnine_unit ninexnine_unit_2445(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10029)
);

ninexnine_unit ninexnine_unit_2446(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11029)
);

ninexnine_unit ninexnine_unit_2447(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12029)
);

assign C1029=c10029+c11029+c12029;
assign A1029=(C1029>=0)?1:0;

assign P2029=A1029;

ninexnine_unit ninexnine_unit_2448(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10039)
);

ninexnine_unit ninexnine_unit_2449(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11039)
);

ninexnine_unit ninexnine_unit_2450(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12039)
);

assign C1039=c10039+c11039+c12039;
assign A1039=(C1039>=0)?1:0;

assign P2039=A1039;

ninexnine_unit ninexnine_unit_2451(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10049)
);

ninexnine_unit ninexnine_unit_2452(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11049)
);

ninexnine_unit ninexnine_unit_2453(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12049)
);

assign C1049=c10049+c11049+c12049;
assign A1049=(C1049>=0)?1:0;

assign P2049=A1049;

ninexnine_unit ninexnine_unit_2454(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10109)
);

ninexnine_unit ninexnine_unit_2455(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11109)
);

ninexnine_unit ninexnine_unit_2456(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12109)
);

assign C1109=c10109+c11109+c12109;
assign A1109=(C1109>=0)?1:0;

assign P2109=A1109;

ninexnine_unit ninexnine_unit_2457(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10119)
);

ninexnine_unit ninexnine_unit_2458(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11119)
);

ninexnine_unit ninexnine_unit_2459(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12119)
);

assign C1119=c10119+c11119+c12119;
assign A1119=(C1119>=0)?1:0;

assign P2119=A1119;

ninexnine_unit ninexnine_unit_2460(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10129)
);

ninexnine_unit ninexnine_unit_2461(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11129)
);

ninexnine_unit ninexnine_unit_2462(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12129)
);

assign C1129=c10129+c11129+c12129;
assign A1129=(C1129>=0)?1:0;

assign P2129=A1129;

ninexnine_unit ninexnine_unit_2463(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10139)
);

ninexnine_unit ninexnine_unit_2464(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11139)
);

ninexnine_unit ninexnine_unit_2465(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12139)
);

assign C1139=c10139+c11139+c12139;
assign A1139=(C1139>=0)?1:0;

assign P2139=A1139;

ninexnine_unit ninexnine_unit_2466(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10149)
);

ninexnine_unit ninexnine_unit_2467(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11149)
);

ninexnine_unit ninexnine_unit_2468(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12149)
);

assign C1149=c10149+c11149+c12149;
assign A1149=(C1149>=0)?1:0;

assign P2149=A1149;

ninexnine_unit ninexnine_unit_2469(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10209)
);

ninexnine_unit ninexnine_unit_2470(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11209)
);

ninexnine_unit ninexnine_unit_2471(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12209)
);

assign C1209=c10209+c11209+c12209;
assign A1209=(C1209>=0)?1:0;

assign P2209=A1209;

ninexnine_unit ninexnine_unit_2472(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10219)
);

ninexnine_unit ninexnine_unit_2473(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11219)
);

ninexnine_unit ninexnine_unit_2474(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12219)
);

assign C1219=c10219+c11219+c12219;
assign A1219=(C1219>=0)?1:0;

assign P2219=A1219;

ninexnine_unit ninexnine_unit_2475(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10229)
);

ninexnine_unit ninexnine_unit_2476(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11229)
);

ninexnine_unit ninexnine_unit_2477(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12229)
);

assign C1229=c10229+c11229+c12229;
assign A1229=(C1229>=0)?1:0;

assign P2229=A1229;

ninexnine_unit ninexnine_unit_2478(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10239)
);

ninexnine_unit ninexnine_unit_2479(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11239)
);

ninexnine_unit ninexnine_unit_2480(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12239)
);

assign C1239=c10239+c11239+c12239;
assign A1239=(C1239>=0)?1:0;

assign P2239=A1239;

ninexnine_unit ninexnine_unit_2481(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10249)
);

ninexnine_unit ninexnine_unit_2482(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11249)
);

ninexnine_unit ninexnine_unit_2483(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12249)
);

assign C1249=c10249+c11249+c12249;
assign A1249=(C1249>=0)?1:0;

assign P2249=A1249;

ninexnine_unit ninexnine_unit_2484(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10309)
);

ninexnine_unit ninexnine_unit_2485(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11309)
);

ninexnine_unit ninexnine_unit_2486(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12309)
);

assign C1309=c10309+c11309+c12309;
assign A1309=(C1309>=0)?1:0;

assign P2309=A1309;

ninexnine_unit ninexnine_unit_2487(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10319)
);

ninexnine_unit ninexnine_unit_2488(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11319)
);

ninexnine_unit ninexnine_unit_2489(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12319)
);

assign C1319=c10319+c11319+c12319;
assign A1319=(C1319>=0)?1:0;

assign P2319=A1319;

ninexnine_unit ninexnine_unit_2490(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10329)
);

ninexnine_unit ninexnine_unit_2491(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11329)
);

ninexnine_unit ninexnine_unit_2492(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12329)
);

assign C1329=c10329+c11329+c12329;
assign A1329=(C1329>=0)?1:0;

assign P2329=A1329;

ninexnine_unit ninexnine_unit_2493(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10339)
);

ninexnine_unit ninexnine_unit_2494(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11339)
);

ninexnine_unit ninexnine_unit_2495(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12339)
);

assign C1339=c10339+c11339+c12339;
assign A1339=(C1339>=0)?1:0;

assign P2339=A1339;

ninexnine_unit ninexnine_unit_2496(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10349)
);

ninexnine_unit ninexnine_unit_2497(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11349)
);

ninexnine_unit ninexnine_unit_2498(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12349)
);

assign C1349=c10349+c11349+c12349;
assign A1349=(C1349>=0)?1:0;

assign P2349=A1349;

ninexnine_unit ninexnine_unit_2499(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10409)
);

ninexnine_unit ninexnine_unit_2500(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11409)
);

ninexnine_unit ninexnine_unit_2501(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12409)
);

assign C1409=c10409+c11409+c12409;
assign A1409=(C1409>=0)?1:0;

assign P2409=A1409;

ninexnine_unit ninexnine_unit_2502(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10419)
);

ninexnine_unit ninexnine_unit_2503(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11419)
);

ninexnine_unit ninexnine_unit_2504(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12419)
);

assign C1419=c10419+c11419+c12419;
assign A1419=(C1419>=0)?1:0;

assign P2419=A1419;

ninexnine_unit ninexnine_unit_2505(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10429)
);

ninexnine_unit ninexnine_unit_2506(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11429)
);

ninexnine_unit ninexnine_unit_2507(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12429)
);

assign C1429=c10429+c11429+c12429;
assign A1429=(C1429>=0)?1:0;

assign P2429=A1429;

ninexnine_unit ninexnine_unit_2508(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10439)
);

ninexnine_unit ninexnine_unit_2509(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11439)
);

ninexnine_unit ninexnine_unit_2510(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12439)
);

assign C1439=c10439+c11439+c12439;
assign A1439=(C1439>=0)?1:0;

assign P2439=A1439;

ninexnine_unit ninexnine_unit_2511(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W19000),
				.b1(W19010),
				.b2(W19020),
				.b3(W19100),
				.b4(W19110),
				.b5(W19120),
				.b6(W19200),
				.b7(W19210),
				.b8(W19220),
				.c(c10449)
);

ninexnine_unit ninexnine_unit_2512(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W19001),
				.b1(W19011),
				.b2(W19021),
				.b3(W19101),
				.b4(W19111),
				.b5(W19121),
				.b6(W19201),
				.b7(W19211),
				.b8(W19221),
				.c(c11449)
);

ninexnine_unit ninexnine_unit_2513(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W19002),
				.b1(W19012),
				.b2(W19022),
				.b3(W19102),
				.b4(W19112),
				.b5(W19122),
				.b6(W19202),
				.b7(W19212),
				.b8(W19222),
				.c(c12449)
);

assign C1449=c10449+c11449+c12449;
assign A1449=(C1449>=0)?1:0;

assign P2449=A1449;

ninexnine_unit ninexnine_unit_2514(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1000A)
);

ninexnine_unit ninexnine_unit_2515(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1100A)
);

ninexnine_unit ninexnine_unit_2516(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1200A)
);

assign C100A=c1000A+c1100A+c1200A;
assign A100A=(C100A>=0)?1:0;

assign P200A=A100A;

ninexnine_unit ninexnine_unit_2517(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1001A)
);

ninexnine_unit ninexnine_unit_2518(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1101A)
);

ninexnine_unit ninexnine_unit_2519(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1201A)
);

assign C101A=c1001A+c1101A+c1201A;
assign A101A=(C101A>=0)?1:0;

assign P201A=A101A;

ninexnine_unit ninexnine_unit_2520(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1002A)
);

ninexnine_unit ninexnine_unit_2521(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1102A)
);

ninexnine_unit ninexnine_unit_2522(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1202A)
);

assign C102A=c1002A+c1102A+c1202A;
assign A102A=(C102A>=0)?1:0;

assign P202A=A102A;

ninexnine_unit ninexnine_unit_2523(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1003A)
);

ninexnine_unit ninexnine_unit_2524(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1103A)
);

ninexnine_unit ninexnine_unit_2525(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1203A)
);

assign C103A=c1003A+c1103A+c1203A;
assign A103A=(C103A>=0)?1:0;

assign P203A=A103A;

ninexnine_unit ninexnine_unit_2526(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1004A)
);

ninexnine_unit ninexnine_unit_2527(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1104A)
);

ninexnine_unit ninexnine_unit_2528(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1204A)
);

assign C104A=c1004A+c1104A+c1204A;
assign A104A=(C104A>=0)?1:0;

assign P204A=A104A;

ninexnine_unit ninexnine_unit_2529(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1010A)
);

ninexnine_unit ninexnine_unit_2530(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1110A)
);

ninexnine_unit ninexnine_unit_2531(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1210A)
);

assign C110A=c1010A+c1110A+c1210A;
assign A110A=(C110A>=0)?1:0;

assign P210A=A110A;

ninexnine_unit ninexnine_unit_2532(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1011A)
);

ninexnine_unit ninexnine_unit_2533(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1111A)
);

ninexnine_unit ninexnine_unit_2534(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1211A)
);

assign C111A=c1011A+c1111A+c1211A;
assign A111A=(C111A>=0)?1:0;

assign P211A=A111A;

ninexnine_unit ninexnine_unit_2535(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1012A)
);

ninexnine_unit ninexnine_unit_2536(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1112A)
);

ninexnine_unit ninexnine_unit_2537(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1212A)
);

assign C112A=c1012A+c1112A+c1212A;
assign A112A=(C112A>=0)?1:0;

assign P212A=A112A;

ninexnine_unit ninexnine_unit_2538(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1013A)
);

ninexnine_unit ninexnine_unit_2539(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1113A)
);

ninexnine_unit ninexnine_unit_2540(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1213A)
);

assign C113A=c1013A+c1113A+c1213A;
assign A113A=(C113A>=0)?1:0;

assign P213A=A113A;

ninexnine_unit ninexnine_unit_2541(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1014A)
);

ninexnine_unit ninexnine_unit_2542(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1114A)
);

ninexnine_unit ninexnine_unit_2543(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1214A)
);

assign C114A=c1014A+c1114A+c1214A;
assign A114A=(C114A>=0)?1:0;

assign P214A=A114A;

ninexnine_unit ninexnine_unit_2544(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1020A)
);

ninexnine_unit ninexnine_unit_2545(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1120A)
);

ninexnine_unit ninexnine_unit_2546(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1220A)
);

assign C120A=c1020A+c1120A+c1220A;
assign A120A=(C120A>=0)?1:0;

assign P220A=A120A;

ninexnine_unit ninexnine_unit_2547(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1021A)
);

ninexnine_unit ninexnine_unit_2548(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1121A)
);

ninexnine_unit ninexnine_unit_2549(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1221A)
);

assign C121A=c1021A+c1121A+c1221A;
assign A121A=(C121A>=0)?1:0;

assign P221A=A121A;

ninexnine_unit ninexnine_unit_2550(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1022A)
);

ninexnine_unit ninexnine_unit_2551(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1122A)
);

ninexnine_unit ninexnine_unit_2552(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1222A)
);

assign C122A=c1022A+c1122A+c1222A;
assign A122A=(C122A>=0)?1:0;

assign P222A=A122A;

ninexnine_unit ninexnine_unit_2553(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1023A)
);

ninexnine_unit ninexnine_unit_2554(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1123A)
);

ninexnine_unit ninexnine_unit_2555(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1223A)
);

assign C123A=c1023A+c1123A+c1223A;
assign A123A=(C123A>=0)?1:0;

assign P223A=A123A;

ninexnine_unit ninexnine_unit_2556(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1024A)
);

ninexnine_unit ninexnine_unit_2557(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1124A)
);

ninexnine_unit ninexnine_unit_2558(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1224A)
);

assign C124A=c1024A+c1124A+c1224A;
assign A124A=(C124A>=0)?1:0;

assign P224A=A124A;

ninexnine_unit ninexnine_unit_2559(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1030A)
);

ninexnine_unit ninexnine_unit_2560(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1130A)
);

ninexnine_unit ninexnine_unit_2561(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1230A)
);

assign C130A=c1030A+c1130A+c1230A;
assign A130A=(C130A>=0)?1:0;

assign P230A=A130A;

ninexnine_unit ninexnine_unit_2562(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1031A)
);

ninexnine_unit ninexnine_unit_2563(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1131A)
);

ninexnine_unit ninexnine_unit_2564(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1231A)
);

assign C131A=c1031A+c1131A+c1231A;
assign A131A=(C131A>=0)?1:0;

assign P231A=A131A;

ninexnine_unit ninexnine_unit_2565(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1032A)
);

ninexnine_unit ninexnine_unit_2566(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1132A)
);

ninexnine_unit ninexnine_unit_2567(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1232A)
);

assign C132A=c1032A+c1132A+c1232A;
assign A132A=(C132A>=0)?1:0;

assign P232A=A132A;

ninexnine_unit ninexnine_unit_2568(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1033A)
);

ninexnine_unit ninexnine_unit_2569(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1133A)
);

ninexnine_unit ninexnine_unit_2570(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1233A)
);

assign C133A=c1033A+c1133A+c1233A;
assign A133A=(C133A>=0)?1:0;

assign P233A=A133A;

ninexnine_unit ninexnine_unit_2571(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1034A)
);

ninexnine_unit ninexnine_unit_2572(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1134A)
);

ninexnine_unit ninexnine_unit_2573(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1234A)
);

assign C134A=c1034A+c1134A+c1234A;
assign A134A=(C134A>=0)?1:0;

assign P234A=A134A;

ninexnine_unit ninexnine_unit_2574(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1040A)
);

ninexnine_unit ninexnine_unit_2575(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1140A)
);

ninexnine_unit ninexnine_unit_2576(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1240A)
);

assign C140A=c1040A+c1140A+c1240A;
assign A140A=(C140A>=0)?1:0;

assign P240A=A140A;

ninexnine_unit ninexnine_unit_2577(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1041A)
);

ninexnine_unit ninexnine_unit_2578(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1141A)
);

ninexnine_unit ninexnine_unit_2579(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1241A)
);

assign C141A=c1041A+c1141A+c1241A;
assign A141A=(C141A>=0)?1:0;

assign P241A=A141A;

ninexnine_unit ninexnine_unit_2580(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1042A)
);

ninexnine_unit ninexnine_unit_2581(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1142A)
);

ninexnine_unit ninexnine_unit_2582(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1242A)
);

assign C142A=c1042A+c1142A+c1242A;
assign A142A=(C142A>=0)?1:0;

assign P242A=A142A;

ninexnine_unit ninexnine_unit_2583(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1043A)
);

ninexnine_unit ninexnine_unit_2584(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1143A)
);

ninexnine_unit ninexnine_unit_2585(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1243A)
);

assign C143A=c1043A+c1143A+c1243A;
assign A143A=(C143A>=0)?1:0;

assign P243A=A143A;

ninexnine_unit ninexnine_unit_2586(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W1A000),
				.b1(W1A010),
				.b2(W1A020),
				.b3(W1A100),
				.b4(W1A110),
				.b5(W1A120),
				.b6(W1A200),
				.b7(W1A210),
				.b8(W1A220),
				.c(c1044A)
);

ninexnine_unit ninexnine_unit_2587(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W1A001),
				.b1(W1A011),
				.b2(W1A021),
				.b3(W1A101),
				.b4(W1A111),
				.b5(W1A121),
				.b6(W1A201),
				.b7(W1A211),
				.b8(W1A221),
				.c(c1144A)
);

ninexnine_unit ninexnine_unit_2588(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W1A002),
				.b1(W1A012),
				.b2(W1A022),
				.b3(W1A102),
				.b4(W1A112),
				.b5(W1A122),
				.b6(W1A202),
				.b7(W1A212),
				.b8(W1A222),
				.c(c1244A)
);

assign C144A=c1044A+c1144A+c1244A;
assign A144A=(C144A>=0)?1:0;

assign P244A=A144A;

ninexnine_unit ninexnine_unit_2589(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1000B)
);

ninexnine_unit ninexnine_unit_2590(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1100B)
);

ninexnine_unit ninexnine_unit_2591(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1200B)
);

assign C100B=c1000B+c1100B+c1200B;
assign A100B=(C100B>=0)?1:0;

assign P200B=A100B;

ninexnine_unit ninexnine_unit_2592(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1001B)
);

ninexnine_unit ninexnine_unit_2593(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1101B)
);

ninexnine_unit ninexnine_unit_2594(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1201B)
);

assign C101B=c1001B+c1101B+c1201B;
assign A101B=(C101B>=0)?1:0;

assign P201B=A101B;

ninexnine_unit ninexnine_unit_2595(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1002B)
);

ninexnine_unit ninexnine_unit_2596(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1102B)
);

ninexnine_unit ninexnine_unit_2597(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1202B)
);

assign C102B=c1002B+c1102B+c1202B;
assign A102B=(C102B>=0)?1:0;

assign P202B=A102B;

ninexnine_unit ninexnine_unit_2598(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1003B)
);

ninexnine_unit ninexnine_unit_2599(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1103B)
);

ninexnine_unit ninexnine_unit_2600(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1203B)
);

assign C103B=c1003B+c1103B+c1203B;
assign A103B=(C103B>=0)?1:0;

assign P203B=A103B;

ninexnine_unit ninexnine_unit_2601(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1004B)
);

ninexnine_unit ninexnine_unit_2602(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1104B)
);

ninexnine_unit ninexnine_unit_2603(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1204B)
);

assign C104B=c1004B+c1104B+c1204B;
assign A104B=(C104B>=0)?1:0;

assign P204B=A104B;

ninexnine_unit ninexnine_unit_2604(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1010B)
);

ninexnine_unit ninexnine_unit_2605(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1110B)
);

ninexnine_unit ninexnine_unit_2606(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1210B)
);

assign C110B=c1010B+c1110B+c1210B;
assign A110B=(C110B>=0)?1:0;

assign P210B=A110B;

ninexnine_unit ninexnine_unit_2607(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1011B)
);

ninexnine_unit ninexnine_unit_2608(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1111B)
);

ninexnine_unit ninexnine_unit_2609(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1211B)
);

assign C111B=c1011B+c1111B+c1211B;
assign A111B=(C111B>=0)?1:0;

assign P211B=A111B;

ninexnine_unit ninexnine_unit_2610(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1012B)
);

ninexnine_unit ninexnine_unit_2611(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1112B)
);

ninexnine_unit ninexnine_unit_2612(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1212B)
);

assign C112B=c1012B+c1112B+c1212B;
assign A112B=(C112B>=0)?1:0;

assign P212B=A112B;

ninexnine_unit ninexnine_unit_2613(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1013B)
);

ninexnine_unit ninexnine_unit_2614(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1113B)
);

ninexnine_unit ninexnine_unit_2615(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1213B)
);

assign C113B=c1013B+c1113B+c1213B;
assign A113B=(C113B>=0)?1:0;

assign P213B=A113B;

ninexnine_unit ninexnine_unit_2616(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1014B)
);

ninexnine_unit ninexnine_unit_2617(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1114B)
);

ninexnine_unit ninexnine_unit_2618(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1214B)
);

assign C114B=c1014B+c1114B+c1214B;
assign A114B=(C114B>=0)?1:0;

assign P214B=A114B;

ninexnine_unit ninexnine_unit_2619(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1020B)
);

ninexnine_unit ninexnine_unit_2620(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1120B)
);

ninexnine_unit ninexnine_unit_2621(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1220B)
);

assign C120B=c1020B+c1120B+c1220B;
assign A120B=(C120B>=0)?1:0;

assign P220B=A120B;

ninexnine_unit ninexnine_unit_2622(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1021B)
);

ninexnine_unit ninexnine_unit_2623(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1121B)
);

ninexnine_unit ninexnine_unit_2624(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1221B)
);

assign C121B=c1021B+c1121B+c1221B;
assign A121B=(C121B>=0)?1:0;

assign P221B=A121B;

ninexnine_unit ninexnine_unit_2625(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1022B)
);

ninexnine_unit ninexnine_unit_2626(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1122B)
);

ninexnine_unit ninexnine_unit_2627(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1222B)
);

assign C122B=c1022B+c1122B+c1222B;
assign A122B=(C122B>=0)?1:0;

assign P222B=A122B;

ninexnine_unit ninexnine_unit_2628(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1023B)
);

ninexnine_unit ninexnine_unit_2629(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1123B)
);

ninexnine_unit ninexnine_unit_2630(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1223B)
);

assign C123B=c1023B+c1123B+c1223B;
assign A123B=(C123B>=0)?1:0;

assign P223B=A123B;

ninexnine_unit ninexnine_unit_2631(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1024B)
);

ninexnine_unit ninexnine_unit_2632(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1124B)
);

ninexnine_unit ninexnine_unit_2633(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1224B)
);

assign C124B=c1024B+c1124B+c1224B;
assign A124B=(C124B>=0)?1:0;

assign P224B=A124B;

ninexnine_unit ninexnine_unit_2634(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1030B)
);

ninexnine_unit ninexnine_unit_2635(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1130B)
);

ninexnine_unit ninexnine_unit_2636(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1230B)
);

assign C130B=c1030B+c1130B+c1230B;
assign A130B=(C130B>=0)?1:0;

assign P230B=A130B;

ninexnine_unit ninexnine_unit_2637(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1031B)
);

ninexnine_unit ninexnine_unit_2638(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1131B)
);

ninexnine_unit ninexnine_unit_2639(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1231B)
);

assign C131B=c1031B+c1131B+c1231B;
assign A131B=(C131B>=0)?1:0;

assign P231B=A131B;

ninexnine_unit ninexnine_unit_2640(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1032B)
);

ninexnine_unit ninexnine_unit_2641(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1132B)
);

ninexnine_unit ninexnine_unit_2642(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1232B)
);

assign C132B=c1032B+c1132B+c1232B;
assign A132B=(C132B>=0)?1:0;

assign P232B=A132B;

ninexnine_unit ninexnine_unit_2643(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1033B)
);

ninexnine_unit ninexnine_unit_2644(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1133B)
);

ninexnine_unit ninexnine_unit_2645(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1233B)
);

assign C133B=c1033B+c1133B+c1233B;
assign A133B=(C133B>=0)?1:0;

assign P233B=A133B;

ninexnine_unit ninexnine_unit_2646(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1034B)
);

ninexnine_unit ninexnine_unit_2647(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1134B)
);

ninexnine_unit ninexnine_unit_2648(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1234B)
);

assign C134B=c1034B+c1134B+c1234B;
assign A134B=(C134B>=0)?1:0;

assign P234B=A134B;

ninexnine_unit ninexnine_unit_2649(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1040B)
);

ninexnine_unit ninexnine_unit_2650(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1140B)
);

ninexnine_unit ninexnine_unit_2651(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1240B)
);

assign C140B=c1040B+c1140B+c1240B;
assign A140B=(C140B>=0)?1:0;

assign P240B=A140B;

ninexnine_unit ninexnine_unit_2652(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1041B)
);

ninexnine_unit ninexnine_unit_2653(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1141B)
);

ninexnine_unit ninexnine_unit_2654(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1241B)
);

assign C141B=c1041B+c1141B+c1241B;
assign A141B=(C141B>=0)?1:0;

assign P241B=A141B;

ninexnine_unit ninexnine_unit_2655(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1042B)
);

ninexnine_unit ninexnine_unit_2656(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1142B)
);

ninexnine_unit ninexnine_unit_2657(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1242B)
);

assign C142B=c1042B+c1142B+c1242B;
assign A142B=(C142B>=0)?1:0;

assign P242B=A142B;

ninexnine_unit ninexnine_unit_2658(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1043B)
);

ninexnine_unit ninexnine_unit_2659(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1143B)
);

ninexnine_unit ninexnine_unit_2660(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1243B)
);

assign C143B=c1043B+c1143B+c1243B;
assign A143B=(C143B>=0)?1:0;

assign P243B=A143B;

ninexnine_unit ninexnine_unit_2661(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W1B000),
				.b1(W1B010),
				.b2(W1B020),
				.b3(W1B100),
				.b4(W1B110),
				.b5(W1B120),
				.b6(W1B200),
				.b7(W1B210),
				.b8(W1B220),
				.c(c1044B)
);

ninexnine_unit ninexnine_unit_2662(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W1B001),
				.b1(W1B011),
				.b2(W1B021),
				.b3(W1B101),
				.b4(W1B111),
				.b5(W1B121),
				.b6(W1B201),
				.b7(W1B211),
				.b8(W1B221),
				.c(c1144B)
);

ninexnine_unit ninexnine_unit_2663(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W1B002),
				.b1(W1B012),
				.b2(W1B022),
				.b3(W1B102),
				.b4(W1B112),
				.b5(W1B122),
				.b6(W1B202),
				.b7(W1B212),
				.b8(W1B222),
				.c(c1244B)
);

assign C144B=c1044B+c1144B+c1244B;
assign A144B=(C144B>=0)?1:0;

assign P244B=A144B;

ninexnine_unit ninexnine_unit_2664(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1000C)
);

ninexnine_unit ninexnine_unit_2665(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1100C)
);

ninexnine_unit ninexnine_unit_2666(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1200C)
);

assign C100C=c1000C+c1100C+c1200C;
assign A100C=(C100C>=0)?1:0;

assign P200C=A100C;

ninexnine_unit ninexnine_unit_2667(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1001C)
);

ninexnine_unit ninexnine_unit_2668(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1101C)
);

ninexnine_unit ninexnine_unit_2669(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1201C)
);

assign C101C=c1001C+c1101C+c1201C;
assign A101C=(C101C>=0)?1:0;

assign P201C=A101C;

ninexnine_unit ninexnine_unit_2670(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1002C)
);

ninexnine_unit ninexnine_unit_2671(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1102C)
);

ninexnine_unit ninexnine_unit_2672(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1202C)
);

assign C102C=c1002C+c1102C+c1202C;
assign A102C=(C102C>=0)?1:0;

assign P202C=A102C;

ninexnine_unit ninexnine_unit_2673(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1003C)
);

ninexnine_unit ninexnine_unit_2674(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1103C)
);

ninexnine_unit ninexnine_unit_2675(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1203C)
);

assign C103C=c1003C+c1103C+c1203C;
assign A103C=(C103C>=0)?1:0;

assign P203C=A103C;

ninexnine_unit ninexnine_unit_2676(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1004C)
);

ninexnine_unit ninexnine_unit_2677(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1104C)
);

ninexnine_unit ninexnine_unit_2678(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1204C)
);

assign C104C=c1004C+c1104C+c1204C;
assign A104C=(C104C>=0)?1:0;

assign P204C=A104C;

ninexnine_unit ninexnine_unit_2679(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1010C)
);

ninexnine_unit ninexnine_unit_2680(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1110C)
);

ninexnine_unit ninexnine_unit_2681(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1210C)
);

assign C110C=c1010C+c1110C+c1210C;
assign A110C=(C110C>=0)?1:0;

assign P210C=A110C;

ninexnine_unit ninexnine_unit_2682(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1011C)
);

ninexnine_unit ninexnine_unit_2683(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1111C)
);

ninexnine_unit ninexnine_unit_2684(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1211C)
);

assign C111C=c1011C+c1111C+c1211C;
assign A111C=(C111C>=0)?1:0;

assign P211C=A111C;

ninexnine_unit ninexnine_unit_2685(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1012C)
);

ninexnine_unit ninexnine_unit_2686(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1112C)
);

ninexnine_unit ninexnine_unit_2687(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1212C)
);

assign C112C=c1012C+c1112C+c1212C;
assign A112C=(C112C>=0)?1:0;

assign P212C=A112C;

ninexnine_unit ninexnine_unit_2688(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1013C)
);

ninexnine_unit ninexnine_unit_2689(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1113C)
);

ninexnine_unit ninexnine_unit_2690(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1213C)
);

assign C113C=c1013C+c1113C+c1213C;
assign A113C=(C113C>=0)?1:0;

assign P213C=A113C;

ninexnine_unit ninexnine_unit_2691(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1014C)
);

ninexnine_unit ninexnine_unit_2692(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1114C)
);

ninexnine_unit ninexnine_unit_2693(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1214C)
);

assign C114C=c1014C+c1114C+c1214C;
assign A114C=(C114C>=0)?1:0;

assign P214C=A114C;

ninexnine_unit ninexnine_unit_2694(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1020C)
);

ninexnine_unit ninexnine_unit_2695(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1120C)
);

ninexnine_unit ninexnine_unit_2696(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1220C)
);

assign C120C=c1020C+c1120C+c1220C;
assign A120C=(C120C>=0)?1:0;

assign P220C=A120C;

ninexnine_unit ninexnine_unit_2697(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1021C)
);

ninexnine_unit ninexnine_unit_2698(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1121C)
);

ninexnine_unit ninexnine_unit_2699(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1221C)
);

assign C121C=c1021C+c1121C+c1221C;
assign A121C=(C121C>=0)?1:0;

assign P221C=A121C;

ninexnine_unit ninexnine_unit_2700(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1022C)
);

ninexnine_unit ninexnine_unit_2701(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1122C)
);

ninexnine_unit ninexnine_unit_2702(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1222C)
);

assign C122C=c1022C+c1122C+c1222C;
assign A122C=(C122C>=0)?1:0;

assign P222C=A122C;

ninexnine_unit ninexnine_unit_2703(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1023C)
);

ninexnine_unit ninexnine_unit_2704(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1123C)
);

ninexnine_unit ninexnine_unit_2705(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1223C)
);

assign C123C=c1023C+c1123C+c1223C;
assign A123C=(C123C>=0)?1:0;

assign P223C=A123C;

ninexnine_unit ninexnine_unit_2706(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1024C)
);

ninexnine_unit ninexnine_unit_2707(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1124C)
);

ninexnine_unit ninexnine_unit_2708(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1224C)
);

assign C124C=c1024C+c1124C+c1224C;
assign A124C=(C124C>=0)?1:0;

assign P224C=A124C;

ninexnine_unit ninexnine_unit_2709(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1030C)
);

ninexnine_unit ninexnine_unit_2710(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1130C)
);

ninexnine_unit ninexnine_unit_2711(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1230C)
);

assign C130C=c1030C+c1130C+c1230C;
assign A130C=(C130C>=0)?1:0;

assign P230C=A130C;

ninexnine_unit ninexnine_unit_2712(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1031C)
);

ninexnine_unit ninexnine_unit_2713(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1131C)
);

ninexnine_unit ninexnine_unit_2714(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1231C)
);

assign C131C=c1031C+c1131C+c1231C;
assign A131C=(C131C>=0)?1:0;

assign P231C=A131C;

ninexnine_unit ninexnine_unit_2715(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1032C)
);

ninexnine_unit ninexnine_unit_2716(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1132C)
);

ninexnine_unit ninexnine_unit_2717(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1232C)
);

assign C132C=c1032C+c1132C+c1232C;
assign A132C=(C132C>=0)?1:0;

assign P232C=A132C;

ninexnine_unit ninexnine_unit_2718(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1033C)
);

ninexnine_unit ninexnine_unit_2719(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1133C)
);

ninexnine_unit ninexnine_unit_2720(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1233C)
);

assign C133C=c1033C+c1133C+c1233C;
assign A133C=(C133C>=0)?1:0;

assign P233C=A133C;

ninexnine_unit ninexnine_unit_2721(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1034C)
);

ninexnine_unit ninexnine_unit_2722(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1134C)
);

ninexnine_unit ninexnine_unit_2723(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1234C)
);

assign C134C=c1034C+c1134C+c1234C;
assign A134C=(C134C>=0)?1:0;

assign P234C=A134C;

ninexnine_unit ninexnine_unit_2724(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1040C)
);

ninexnine_unit ninexnine_unit_2725(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1140C)
);

ninexnine_unit ninexnine_unit_2726(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1240C)
);

assign C140C=c1040C+c1140C+c1240C;
assign A140C=(C140C>=0)?1:0;

assign P240C=A140C;

ninexnine_unit ninexnine_unit_2727(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1041C)
);

ninexnine_unit ninexnine_unit_2728(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1141C)
);

ninexnine_unit ninexnine_unit_2729(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1241C)
);

assign C141C=c1041C+c1141C+c1241C;
assign A141C=(C141C>=0)?1:0;

assign P241C=A141C;

ninexnine_unit ninexnine_unit_2730(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1042C)
);

ninexnine_unit ninexnine_unit_2731(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1142C)
);

ninexnine_unit ninexnine_unit_2732(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1242C)
);

assign C142C=c1042C+c1142C+c1242C;
assign A142C=(C142C>=0)?1:0;

assign P242C=A142C;

ninexnine_unit ninexnine_unit_2733(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1043C)
);

ninexnine_unit ninexnine_unit_2734(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1143C)
);

ninexnine_unit ninexnine_unit_2735(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1243C)
);

assign C143C=c1043C+c1143C+c1243C;
assign A143C=(C143C>=0)?1:0;

assign P243C=A143C;

ninexnine_unit ninexnine_unit_2736(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W1C000),
				.b1(W1C010),
				.b2(W1C020),
				.b3(W1C100),
				.b4(W1C110),
				.b5(W1C120),
				.b6(W1C200),
				.b7(W1C210),
				.b8(W1C220),
				.c(c1044C)
);

ninexnine_unit ninexnine_unit_2737(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W1C001),
				.b1(W1C011),
				.b2(W1C021),
				.b3(W1C101),
				.b4(W1C111),
				.b5(W1C121),
				.b6(W1C201),
				.b7(W1C211),
				.b8(W1C221),
				.c(c1144C)
);

ninexnine_unit ninexnine_unit_2738(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W1C002),
				.b1(W1C012),
				.b2(W1C022),
				.b3(W1C102),
				.b4(W1C112),
				.b5(W1C122),
				.b6(W1C202),
				.b7(W1C212),
				.b8(W1C222),
				.c(c1244C)
);

assign C144C=c1044C+c1144C+c1244C;
assign A144C=(C144C>=0)?1:0;

assign P244C=A144C;

ninexnine_unit ninexnine_unit_2739(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1000D)
);

ninexnine_unit ninexnine_unit_2740(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1100D)
);

ninexnine_unit ninexnine_unit_2741(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1200D)
);

assign C100D=c1000D+c1100D+c1200D;
assign A100D=(C100D>=0)?1:0;

assign P200D=A100D;

ninexnine_unit ninexnine_unit_2742(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1001D)
);

ninexnine_unit ninexnine_unit_2743(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1101D)
);

ninexnine_unit ninexnine_unit_2744(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1201D)
);

assign C101D=c1001D+c1101D+c1201D;
assign A101D=(C101D>=0)?1:0;

assign P201D=A101D;

ninexnine_unit ninexnine_unit_2745(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1002D)
);

ninexnine_unit ninexnine_unit_2746(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1102D)
);

ninexnine_unit ninexnine_unit_2747(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1202D)
);

assign C102D=c1002D+c1102D+c1202D;
assign A102D=(C102D>=0)?1:0;

assign P202D=A102D;

ninexnine_unit ninexnine_unit_2748(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1003D)
);

ninexnine_unit ninexnine_unit_2749(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1103D)
);

ninexnine_unit ninexnine_unit_2750(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1203D)
);

assign C103D=c1003D+c1103D+c1203D;
assign A103D=(C103D>=0)?1:0;

assign P203D=A103D;

ninexnine_unit ninexnine_unit_2751(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1004D)
);

ninexnine_unit ninexnine_unit_2752(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1104D)
);

ninexnine_unit ninexnine_unit_2753(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1204D)
);

assign C104D=c1004D+c1104D+c1204D;
assign A104D=(C104D>=0)?1:0;

assign P204D=A104D;

ninexnine_unit ninexnine_unit_2754(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1010D)
);

ninexnine_unit ninexnine_unit_2755(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1110D)
);

ninexnine_unit ninexnine_unit_2756(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1210D)
);

assign C110D=c1010D+c1110D+c1210D;
assign A110D=(C110D>=0)?1:0;

assign P210D=A110D;

ninexnine_unit ninexnine_unit_2757(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1011D)
);

ninexnine_unit ninexnine_unit_2758(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1111D)
);

ninexnine_unit ninexnine_unit_2759(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1211D)
);

assign C111D=c1011D+c1111D+c1211D;
assign A111D=(C111D>=0)?1:0;

assign P211D=A111D;

ninexnine_unit ninexnine_unit_2760(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1012D)
);

ninexnine_unit ninexnine_unit_2761(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1112D)
);

ninexnine_unit ninexnine_unit_2762(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1212D)
);

assign C112D=c1012D+c1112D+c1212D;
assign A112D=(C112D>=0)?1:0;

assign P212D=A112D;

ninexnine_unit ninexnine_unit_2763(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1013D)
);

ninexnine_unit ninexnine_unit_2764(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1113D)
);

ninexnine_unit ninexnine_unit_2765(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1213D)
);

assign C113D=c1013D+c1113D+c1213D;
assign A113D=(C113D>=0)?1:0;

assign P213D=A113D;

ninexnine_unit ninexnine_unit_2766(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1014D)
);

ninexnine_unit ninexnine_unit_2767(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1114D)
);

ninexnine_unit ninexnine_unit_2768(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1214D)
);

assign C114D=c1014D+c1114D+c1214D;
assign A114D=(C114D>=0)?1:0;

assign P214D=A114D;

ninexnine_unit ninexnine_unit_2769(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1020D)
);

ninexnine_unit ninexnine_unit_2770(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1120D)
);

ninexnine_unit ninexnine_unit_2771(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1220D)
);

assign C120D=c1020D+c1120D+c1220D;
assign A120D=(C120D>=0)?1:0;

assign P220D=A120D;

ninexnine_unit ninexnine_unit_2772(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1021D)
);

ninexnine_unit ninexnine_unit_2773(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1121D)
);

ninexnine_unit ninexnine_unit_2774(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1221D)
);

assign C121D=c1021D+c1121D+c1221D;
assign A121D=(C121D>=0)?1:0;

assign P221D=A121D;

ninexnine_unit ninexnine_unit_2775(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1022D)
);

ninexnine_unit ninexnine_unit_2776(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1122D)
);

ninexnine_unit ninexnine_unit_2777(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1222D)
);

assign C122D=c1022D+c1122D+c1222D;
assign A122D=(C122D>=0)?1:0;

assign P222D=A122D;

ninexnine_unit ninexnine_unit_2778(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1023D)
);

ninexnine_unit ninexnine_unit_2779(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1123D)
);

ninexnine_unit ninexnine_unit_2780(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1223D)
);

assign C123D=c1023D+c1123D+c1223D;
assign A123D=(C123D>=0)?1:0;

assign P223D=A123D;

ninexnine_unit ninexnine_unit_2781(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1024D)
);

ninexnine_unit ninexnine_unit_2782(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1124D)
);

ninexnine_unit ninexnine_unit_2783(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1224D)
);

assign C124D=c1024D+c1124D+c1224D;
assign A124D=(C124D>=0)?1:0;

assign P224D=A124D;

ninexnine_unit ninexnine_unit_2784(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1030D)
);

ninexnine_unit ninexnine_unit_2785(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1130D)
);

ninexnine_unit ninexnine_unit_2786(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1230D)
);

assign C130D=c1030D+c1130D+c1230D;
assign A130D=(C130D>=0)?1:0;

assign P230D=A130D;

ninexnine_unit ninexnine_unit_2787(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1031D)
);

ninexnine_unit ninexnine_unit_2788(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1131D)
);

ninexnine_unit ninexnine_unit_2789(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1231D)
);

assign C131D=c1031D+c1131D+c1231D;
assign A131D=(C131D>=0)?1:0;

assign P231D=A131D;

ninexnine_unit ninexnine_unit_2790(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1032D)
);

ninexnine_unit ninexnine_unit_2791(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1132D)
);

ninexnine_unit ninexnine_unit_2792(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1232D)
);

assign C132D=c1032D+c1132D+c1232D;
assign A132D=(C132D>=0)?1:0;

assign P232D=A132D;

ninexnine_unit ninexnine_unit_2793(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1033D)
);

ninexnine_unit ninexnine_unit_2794(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1133D)
);

ninexnine_unit ninexnine_unit_2795(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1233D)
);

assign C133D=c1033D+c1133D+c1233D;
assign A133D=(C133D>=0)?1:0;

assign P233D=A133D;

ninexnine_unit ninexnine_unit_2796(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1034D)
);

ninexnine_unit ninexnine_unit_2797(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1134D)
);

ninexnine_unit ninexnine_unit_2798(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1234D)
);

assign C134D=c1034D+c1134D+c1234D;
assign A134D=(C134D>=0)?1:0;

assign P234D=A134D;

ninexnine_unit ninexnine_unit_2799(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1040D)
);

ninexnine_unit ninexnine_unit_2800(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1140D)
);

ninexnine_unit ninexnine_unit_2801(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1240D)
);

assign C140D=c1040D+c1140D+c1240D;
assign A140D=(C140D>=0)?1:0;

assign P240D=A140D;

ninexnine_unit ninexnine_unit_2802(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1041D)
);

ninexnine_unit ninexnine_unit_2803(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1141D)
);

ninexnine_unit ninexnine_unit_2804(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1241D)
);

assign C141D=c1041D+c1141D+c1241D;
assign A141D=(C141D>=0)?1:0;

assign P241D=A141D;

ninexnine_unit ninexnine_unit_2805(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1042D)
);

ninexnine_unit ninexnine_unit_2806(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1142D)
);

ninexnine_unit ninexnine_unit_2807(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1242D)
);

assign C142D=c1042D+c1142D+c1242D;
assign A142D=(C142D>=0)?1:0;

assign P242D=A142D;

ninexnine_unit ninexnine_unit_2808(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1043D)
);

ninexnine_unit ninexnine_unit_2809(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1143D)
);

ninexnine_unit ninexnine_unit_2810(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1243D)
);

assign C143D=c1043D+c1143D+c1243D;
assign A143D=(C143D>=0)?1:0;

assign P243D=A143D;

ninexnine_unit ninexnine_unit_2811(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W1D000),
				.b1(W1D010),
				.b2(W1D020),
				.b3(W1D100),
				.b4(W1D110),
				.b5(W1D120),
				.b6(W1D200),
				.b7(W1D210),
				.b8(W1D220),
				.c(c1044D)
);

ninexnine_unit ninexnine_unit_2812(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W1D001),
				.b1(W1D011),
				.b2(W1D021),
				.b3(W1D101),
				.b4(W1D111),
				.b5(W1D121),
				.b6(W1D201),
				.b7(W1D211),
				.b8(W1D221),
				.c(c1144D)
);

ninexnine_unit ninexnine_unit_2813(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W1D002),
				.b1(W1D012),
				.b2(W1D022),
				.b3(W1D102),
				.b4(W1D112),
				.b5(W1D122),
				.b6(W1D202),
				.b7(W1D212),
				.b8(W1D222),
				.c(c1244D)
);

assign C144D=c1044D+c1144D+c1244D;
assign A144D=(C144D>=0)?1:0;

assign P244D=A144D;

ninexnine_unit ninexnine_unit_2814(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1000E)
);

ninexnine_unit ninexnine_unit_2815(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1100E)
);

ninexnine_unit ninexnine_unit_2816(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1200E)
);

assign C100E=c1000E+c1100E+c1200E;
assign A100E=(C100E>=0)?1:0;

assign P200E=A100E;

ninexnine_unit ninexnine_unit_2817(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1001E)
);

ninexnine_unit ninexnine_unit_2818(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1101E)
);

ninexnine_unit ninexnine_unit_2819(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1201E)
);

assign C101E=c1001E+c1101E+c1201E;
assign A101E=(C101E>=0)?1:0;

assign P201E=A101E;

ninexnine_unit ninexnine_unit_2820(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1002E)
);

ninexnine_unit ninexnine_unit_2821(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1102E)
);

ninexnine_unit ninexnine_unit_2822(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1202E)
);

assign C102E=c1002E+c1102E+c1202E;
assign A102E=(C102E>=0)?1:0;

assign P202E=A102E;

ninexnine_unit ninexnine_unit_2823(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1003E)
);

ninexnine_unit ninexnine_unit_2824(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1103E)
);

ninexnine_unit ninexnine_unit_2825(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1203E)
);

assign C103E=c1003E+c1103E+c1203E;
assign A103E=(C103E>=0)?1:0;

assign P203E=A103E;

ninexnine_unit ninexnine_unit_2826(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1004E)
);

ninexnine_unit ninexnine_unit_2827(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1104E)
);

ninexnine_unit ninexnine_unit_2828(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1204E)
);

assign C104E=c1004E+c1104E+c1204E;
assign A104E=(C104E>=0)?1:0;

assign P204E=A104E;

ninexnine_unit ninexnine_unit_2829(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1010E)
);

ninexnine_unit ninexnine_unit_2830(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1110E)
);

ninexnine_unit ninexnine_unit_2831(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1210E)
);

assign C110E=c1010E+c1110E+c1210E;
assign A110E=(C110E>=0)?1:0;

assign P210E=A110E;

ninexnine_unit ninexnine_unit_2832(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1011E)
);

ninexnine_unit ninexnine_unit_2833(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1111E)
);

ninexnine_unit ninexnine_unit_2834(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1211E)
);

assign C111E=c1011E+c1111E+c1211E;
assign A111E=(C111E>=0)?1:0;

assign P211E=A111E;

ninexnine_unit ninexnine_unit_2835(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1012E)
);

ninexnine_unit ninexnine_unit_2836(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1112E)
);

ninexnine_unit ninexnine_unit_2837(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1212E)
);

assign C112E=c1012E+c1112E+c1212E;
assign A112E=(C112E>=0)?1:0;

assign P212E=A112E;

ninexnine_unit ninexnine_unit_2838(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1013E)
);

ninexnine_unit ninexnine_unit_2839(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1113E)
);

ninexnine_unit ninexnine_unit_2840(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1213E)
);

assign C113E=c1013E+c1113E+c1213E;
assign A113E=(C113E>=0)?1:0;

assign P213E=A113E;

ninexnine_unit ninexnine_unit_2841(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1014E)
);

ninexnine_unit ninexnine_unit_2842(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1114E)
);

ninexnine_unit ninexnine_unit_2843(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1214E)
);

assign C114E=c1014E+c1114E+c1214E;
assign A114E=(C114E>=0)?1:0;

assign P214E=A114E;

ninexnine_unit ninexnine_unit_2844(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1020E)
);

ninexnine_unit ninexnine_unit_2845(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1120E)
);

ninexnine_unit ninexnine_unit_2846(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1220E)
);

assign C120E=c1020E+c1120E+c1220E;
assign A120E=(C120E>=0)?1:0;

assign P220E=A120E;

ninexnine_unit ninexnine_unit_2847(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1021E)
);

ninexnine_unit ninexnine_unit_2848(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1121E)
);

ninexnine_unit ninexnine_unit_2849(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1221E)
);

assign C121E=c1021E+c1121E+c1221E;
assign A121E=(C121E>=0)?1:0;

assign P221E=A121E;

ninexnine_unit ninexnine_unit_2850(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1022E)
);

ninexnine_unit ninexnine_unit_2851(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1122E)
);

ninexnine_unit ninexnine_unit_2852(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1222E)
);

assign C122E=c1022E+c1122E+c1222E;
assign A122E=(C122E>=0)?1:0;

assign P222E=A122E;

ninexnine_unit ninexnine_unit_2853(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1023E)
);

ninexnine_unit ninexnine_unit_2854(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1123E)
);

ninexnine_unit ninexnine_unit_2855(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1223E)
);

assign C123E=c1023E+c1123E+c1223E;
assign A123E=(C123E>=0)?1:0;

assign P223E=A123E;

ninexnine_unit ninexnine_unit_2856(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1024E)
);

ninexnine_unit ninexnine_unit_2857(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1124E)
);

ninexnine_unit ninexnine_unit_2858(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1224E)
);

assign C124E=c1024E+c1124E+c1224E;
assign A124E=(C124E>=0)?1:0;

assign P224E=A124E;

ninexnine_unit ninexnine_unit_2859(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1030E)
);

ninexnine_unit ninexnine_unit_2860(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1130E)
);

ninexnine_unit ninexnine_unit_2861(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1230E)
);

assign C130E=c1030E+c1130E+c1230E;
assign A130E=(C130E>=0)?1:0;

assign P230E=A130E;

ninexnine_unit ninexnine_unit_2862(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1031E)
);

ninexnine_unit ninexnine_unit_2863(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1131E)
);

ninexnine_unit ninexnine_unit_2864(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1231E)
);

assign C131E=c1031E+c1131E+c1231E;
assign A131E=(C131E>=0)?1:0;

assign P231E=A131E;

ninexnine_unit ninexnine_unit_2865(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1032E)
);

ninexnine_unit ninexnine_unit_2866(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1132E)
);

ninexnine_unit ninexnine_unit_2867(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1232E)
);

assign C132E=c1032E+c1132E+c1232E;
assign A132E=(C132E>=0)?1:0;

assign P232E=A132E;

ninexnine_unit ninexnine_unit_2868(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1033E)
);

ninexnine_unit ninexnine_unit_2869(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1133E)
);

ninexnine_unit ninexnine_unit_2870(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1233E)
);

assign C133E=c1033E+c1133E+c1233E;
assign A133E=(C133E>=0)?1:0;

assign P233E=A133E;

ninexnine_unit ninexnine_unit_2871(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1034E)
);

ninexnine_unit ninexnine_unit_2872(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1134E)
);

ninexnine_unit ninexnine_unit_2873(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1234E)
);

assign C134E=c1034E+c1134E+c1234E;
assign A134E=(C134E>=0)?1:0;

assign P234E=A134E;

ninexnine_unit ninexnine_unit_2874(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1040E)
);

ninexnine_unit ninexnine_unit_2875(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1140E)
);

ninexnine_unit ninexnine_unit_2876(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1240E)
);

assign C140E=c1040E+c1140E+c1240E;
assign A140E=(C140E>=0)?1:0;

assign P240E=A140E;

ninexnine_unit ninexnine_unit_2877(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1041E)
);

ninexnine_unit ninexnine_unit_2878(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1141E)
);

ninexnine_unit ninexnine_unit_2879(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1241E)
);

assign C141E=c1041E+c1141E+c1241E;
assign A141E=(C141E>=0)?1:0;

assign P241E=A141E;

ninexnine_unit ninexnine_unit_2880(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1042E)
);

ninexnine_unit ninexnine_unit_2881(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1142E)
);

ninexnine_unit ninexnine_unit_2882(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1242E)
);

assign C142E=c1042E+c1142E+c1242E;
assign A142E=(C142E>=0)?1:0;

assign P242E=A142E;

ninexnine_unit ninexnine_unit_2883(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1043E)
);

ninexnine_unit ninexnine_unit_2884(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1143E)
);

ninexnine_unit ninexnine_unit_2885(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1243E)
);

assign C143E=c1043E+c1143E+c1243E;
assign A143E=(C143E>=0)?1:0;

assign P243E=A143E;

ninexnine_unit ninexnine_unit_2886(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W1E000),
				.b1(W1E010),
				.b2(W1E020),
				.b3(W1E100),
				.b4(W1E110),
				.b5(W1E120),
				.b6(W1E200),
				.b7(W1E210),
				.b8(W1E220),
				.c(c1044E)
);

ninexnine_unit ninexnine_unit_2887(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W1E001),
				.b1(W1E011),
				.b2(W1E021),
				.b3(W1E101),
				.b4(W1E111),
				.b5(W1E121),
				.b6(W1E201),
				.b7(W1E211),
				.b8(W1E221),
				.c(c1144E)
);

ninexnine_unit ninexnine_unit_2888(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W1E002),
				.b1(W1E012),
				.b2(W1E022),
				.b3(W1E102),
				.b4(W1E112),
				.b5(W1E122),
				.b6(W1E202),
				.b7(W1E212),
				.b8(W1E222),
				.c(c1244E)
);

assign C144E=c1044E+c1144E+c1244E;
assign A144E=(C144E>=0)?1:0;

assign P244E=A144E;

ninexnine_unit ninexnine_unit_2889(
				.clk(clk),
				.rstn(rstn),
				.a0(P1000),
				.a1(P1010),
				.a2(P1020),
				.a3(P1100),
				.a4(P1110),
				.a5(P1120),
				.a6(P1200),
				.a7(P1210),
				.a8(P1220),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1000F)
);

ninexnine_unit ninexnine_unit_2890(
				.clk(clk),
				.rstn(rstn),
				.a0(P1001),
				.a1(P1011),
				.a2(P1021),
				.a3(P1101),
				.a4(P1111),
				.a5(P1121),
				.a6(P1201),
				.a7(P1211),
				.a8(P1221),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1100F)
);

ninexnine_unit ninexnine_unit_2891(
				.clk(clk),
				.rstn(rstn),
				.a0(P1002),
				.a1(P1012),
				.a2(P1022),
				.a3(P1102),
				.a4(P1112),
				.a5(P1122),
				.a6(P1202),
				.a7(P1212),
				.a8(P1222),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1200F)
);

assign C100F=c1000F+c1100F+c1200F;
assign A100F=(C100F>=0)?1:0;

assign P200F=A100F;

ninexnine_unit ninexnine_unit_2892(
				.clk(clk),
				.rstn(rstn),
				.a0(P1010),
				.a1(P1020),
				.a2(P1030),
				.a3(P1110),
				.a4(P1120),
				.a5(P1130),
				.a6(P1210),
				.a7(P1220),
				.a8(P1230),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1001F)
);

ninexnine_unit ninexnine_unit_2893(
				.clk(clk),
				.rstn(rstn),
				.a0(P1011),
				.a1(P1021),
				.a2(P1031),
				.a3(P1111),
				.a4(P1121),
				.a5(P1131),
				.a6(P1211),
				.a7(P1221),
				.a8(P1231),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1101F)
);

ninexnine_unit ninexnine_unit_2894(
				.clk(clk),
				.rstn(rstn),
				.a0(P1012),
				.a1(P1022),
				.a2(P1032),
				.a3(P1112),
				.a4(P1122),
				.a5(P1132),
				.a6(P1212),
				.a7(P1222),
				.a8(P1232),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1201F)
);

assign C101F=c1001F+c1101F+c1201F;
assign A101F=(C101F>=0)?1:0;

assign P201F=A101F;

ninexnine_unit ninexnine_unit_2895(
				.clk(clk),
				.rstn(rstn),
				.a0(P1020),
				.a1(P1030),
				.a2(P1040),
				.a3(P1120),
				.a4(P1130),
				.a5(P1140),
				.a6(P1220),
				.a7(P1230),
				.a8(P1240),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1002F)
);

ninexnine_unit ninexnine_unit_2896(
				.clk(clk),
				.rstn(rstn),
				.a0(P1021),
				.a1(P1031),
				.a2(P1041),
				.a3(P1121),
				.a4(P1131),
				.a5(P1141),
				.a6(P1221),
				.a7(P1231),
				.a8(P1241),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1102F)
);

ninexnine_unit ninexnine_unit_2897(
				.clk(clk),
				.rstn(rstn),
				.a0(P1022),
				.a1(P1032),
				.a2(P1042),
				.a3(P1122),
				.a4(P1132),
				.a5(P1142),
				.a6(P1222),
				.a7(P1232),
				.a8(P1242),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1202F)
);

assign C102F=c1002F+c1102F+c1202F;
assign A102F=(C102F>=0)?1:0;

assign P202F=A102F;

ninexnine_unit ninexnine_unit_2898(
				.clk(clk),
				.rstn(rstn),
				.a0(P1030),
				.a1(P1040),
				.a2(P1050),
				.a3(P1130),
				.a4(P1140),
				.a5(P1150),
				.a6(P1230),
				.a7(P1240),
				.a8(P1250),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1003F)
);

ninexnine_unit ninexnine_unit_2899(
				.clk(clk),
				.rstn(rstn),
				.a0(P1031),
				.a1(P1041),
				.a2(P1051),
				.a3(P1131),
				.a4(P1141),
				.a5(P1151),
				.a6(P1231),
				.a7(P1241),
				.a8(P1251),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1103F)
);

ninexnine_unit ninexnine_unit_2900(
				.clk(clk),
				.rstn(rstn),
				.a0(P1032),
				.a1(P1042),
				.a2(P1052),
				.a3(P1132),
				.a4(P1142),
				.a5(P1152),
				.a6(P1232),
				.a7(P1242),
				.a8(P1252),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1203F)
);

assign C103F=c1003F+c1103F+c1203F;
assign A103F=(C103F>=0)?1:0;

assign P203F=A103F;

ninexnine_unit ninexnine_unit_2901(
				.clk(clk),
				.rstn(rstn),
				.a0(P1040),
				.a1(P1050),
				.a2(P1060),
				.a3(P1140),
				.a4(P1150),
				.a5(P1160),
				.a6(P1240),
				.a7(P1250),
				.a8(P1260),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1004F)
);

ninexnine_unit ninexnine_unit_2902(
				.clk(clk),
				.rstn(rstn),
				.a0(P1041),
				.a1(P1051),
				.a2(P1061),
				.a3(P1141),
				.a4(P1151),
				.a5(P1161),
				.a6(P1241),
				.a7(P1251),
				.a8(P1261),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1104F)
);

ninexnine_unit ninexnine_unit_2903(
				.clk(clk),
				.rstn(rstn),
				.a0(P1042),
				.a1(P1052),
				.a2(P1062),
				.a3(P1142),
				.a4(P1152),
				.a5(P1162),
				.a6(P1242),
				.a7(P1252),
				.a8(P1262),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1204F)
);

assign C104F=c1004F+c1104F+c1204F;
assign A104F=(C104F>=0)?1:0;

assign P204F=A104F;

ninexnine_unit ninexnine_unit_2904(
				.clk(clk),
				.rstn(rstn),
				.a0(P1100),
				.a1(P1110),
				.a2(P1120),
				.a3(P1200),
				.a4(P1210),
				.a5(P1220),
				.a6(P1300),
				.a7(P1310),
				.a8(P1320),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1010F)
);

ninexnine_unit ninexnine_unit_2905(
				.clk(clk),
				.rstn(rstn),
				.a0(P1101),
				.a1(P1111),
				.a2(P1121),
				.a3(P1201),
				.a4(P1211),
				.a5(P1221),
				.a6(P1301),
				.a7(P1311),
				.a8(P1321),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1110F)
);

ninexnine_unit ninexnine_unit_2906(
				.clk(clk),
				.rstn(rstn),
				.a0(P1102),
				.a1(P1112),
				.a2(P1122),
				.a3(P1202),
				.a4(P1212),
				.a5(P1222),
				.a6(P1302),
				.a7(P1312),
				.a8(P1322),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1210F)
);

assign C110F=c1010F+c1110F+c1210F;
assign A110F=(C110F>=0)?1:0;

assign P210F=A110F;

ninexnine_unit ninexnine_unit_2907(
				.clk(clk),
				.rstn(rstn),
				.a0(P1110),
				.a1(P1120),
				.a2(P1130),
				.a3(P1210),
				.a4(P1220),
				.a5(P1230),
				.a6(P1310),
				.a7(P1320),
				.a8(P1330),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1011F)
);

ninexnine_unit ninexnine_unit_2908(
				.clk(clk),
				.rstn(rstn),
				.a0(P1111),
				.a1(P1121),
				.a2(P1131),
				.a3(P1211),
				.a4(P1221),
				.a5(P1231),
				.a6(P1311),
				.a7(P1321),
				.a8(P1331),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1111F)
);

ninexnine_unit ninexnine_unit_2909(
				.clk(clk),
				.rstn(rstn),
				.a0(P1112),
				.a1(P1122),
				.a2(P1132),
				.a3(P1212),
				.a4(P1222),
				.a5(P1232),
				.a6(P1312),
				.a7(P1322),
				.a8(P1332),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1211F)
);

assign C111F=c1011F+c1111F+c1211F;
assign A111F=(C111F>=0)?1:0;

assign P211F=A111F;

ninexnine_unit ninexnine_unit_2910(
				.clk(clk),
				.rstn(rstn),
				.a0(P1120),
				.a1(P1130),
				.a2(P1140),
				.a3(P1220),
				.a4(P1230),
				.a5(P1240),
				.a6(P1320),
				.a7(P1330),
				.a8(P1340),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1012F)
);

ninexnine_unit ninexnine_unit_2911(
				.clk(clk),
				.rstn(rstn),
				.a0(P1121),
				.a1(P1131),
				.a2(P1141),
				.a3(P1221),
				.a4(P1231),
				.a5(P1241),
				.a6(P1321),
				.a7(P1331),
				.a8(P1341),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1112F)
);

ninexnine_unit ninexnine_unit_2912(
				.clk(clk),
				.rstn(rstn),
				.a0(P1122),
				.a1(P1132),
				.a2(P1142),
				.a3(P1222),
				.a4(P1232),
				.a5(P1242),
				.a6(P1322),
				.a7(P1332),
				.a8(P1342),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1212F)
);

assign C112F=c1012F+c1112F+c1212F;
assign A112F=(C112F>=0)?1:0;

assign P212F=A112F;

ninexnine_unit ninexnine_unit_2913(
				.clk(clk),
				.rstn(rstn),
				.a0(P1130),
				.a1(P1140),
				.a2(P1150),
				.a3(P1230),
				.a4(P1240),
				.a5(P1250),
				.a6(P1330),
				.a7(P1340),
				.a8(P1350),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1013F)
);

ninexnine_unit ninexnine_unit_2914(
				.clk(clk),
				.rstn(rstn),
				.a0(P1131),
				.a1(P1141),
				.a2(P1151),
				.a3(P1231),
				.a4(P1241),
				.a5(P1251),
				.a6(P1331),
				.a7(P1341),
				.a8(P1351),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1113F)
);

ninexnine_unit ninexnine_unit_2915(
				.clk(clk),
				.rstn(rstn),
				.a0(P1132),
				.a1(P1142),
				.a2(P1152),
				.a3(P1232),
				.a4(P1242),
				.a5(P1252),
				.a6(P1332),
				.a7(P1342),
				.a8(P1352),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1213F)
);

assign C113F=c1013F+c1113F+c1213F;
assign A113F=(C113F>=0)?1:0;

assign P213F=A113F;

ninexnine_unit ninexnine_unit_2916(
				.clk(clk),
				.rstn(rstn),
				.a0(P1140),
				.a1(P1150),
				.a2(P1160),
				.a3(P1240),
				.a4(P1250),
				.a5(P1260),
				.a6(P1340),
				.a7(P1350),
				.a8(P1360),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1014F)
);

ninexnine_unit ninexnine_unit_2917(
				.clk(clk),
				.rstn(rstn),
				.a0(P1141),
				.a1(P1151),
				.a2(P1161),
				.a3(P1241),
				.a4(P1251),
				.a5(P1261),
				.a6(P1341),
				.a7(P1351),
				.a8(P1361),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1114F)
);

ninexnine_unit ninexnine_unit_2918(
				.clk(clk),
				.rstn(rstn),
				.a0(P1142),
				.a1(P1152),
				.a2(P1162),
				.a3(P1242),
				.a4(P1252),
				.a5(P1262),
				.a6(P1342),
				.a7(P1352),
				.a8(P1362),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1214F)
);

assign C114F=c1014F+c1114F+c1214F;
assign A114F=(C114F>=0)?1:0;

assign P214F=A114F;

ninexnine_unit ninexnine_unit_2919(
				.clk(clk),
				.rstn(rstn),
				.a0(P1200),
				.a1(P1210),
				.a2(P1220),
				.a3(P1300),
				.a4(P1310),
				.a5(P1320),
				.a6(P1400),
				.a7(P1410),
				.a8(P1420),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1020F)
);

ninexnine_unit ninexnine_unit_2920(
				.clk(clk),
				.rstn(rstn),
				.a0(P1201),
				.a1(P1211),
				.a2(P1221),
				.a3(P1301),
				.a4(P1311),
				.a5(P1321),
				.a6(P1401),
				.a7(P1411),
				.a8(P1421),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1120F)
);

ninexnine_unit ninexnine_unit_2921(
				.clk(clk),
				.rstn(rstn),
				.a0(P1202),
				.a1(P1212),
				.a2(P1222),
				.a3(P1302),
				.a4(P1312),
				.a5(P1322),
				.a6(P1402),
				.a7(P1412),
				.a8(P1422),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1220F)
);

assign C120F=c1020F+c1120F+c1220F;
assign A120F=(C120F>=0)?1:0;

assign P220F=A120F;

ninexnine_unit ninexnine_unit_2922(
				.clk(clk),
				.rstn(rstn),
				.a0(P1210),
				.a1(P1220),
				.a2(P1230),
				.a3(P1310),
				.a4(P1320),
				.a5(P1330),
				.a6(P1410),
				.a7(P1420),
				.a8(P1430),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1021F)
);

ninexnine_unit ninexnine_unit_2923(
				.clk(clk),
				.rstn(rstn),
				.a0(P1211),
				.a1(P1221),
				.a2(P1231),
				.a3(P1311),
				.a4(P1321),
				.a5(P1331),
				.a6(P1411),
				.a7(P1421),
				.a8(P1431),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1121F)
);

ninexnine_unit ninexnine_unit_2924(
				.clk(clk),
				.rstn(rstn),
				.a0(P1212),
				.a1(P1222),
				.a2(P1232),
				.a3(P1312),
				.a4(P1322),
				.a5(P1332),
				.a6(P1412),
				.a7(P1422),
				.a8(P1432),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1221F)
);

assign C121F=c1021F+c1121F+c1221F;
assign A121F=(C121F>=0)?1:0;

assign P221F=A121F;

ninexnine_unit ninexnine_unit_2925(
				.clk(clk),
				.rstn(rstn),
				.a0(P1220),
				.a1(P1230),
				.a2(P1240),
				.a3(P1320),
				.a4(P1330),
				.a5(P1340),
				.a6(P1420),
				.a7(P1430),
				.a8(P1440),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1022F)
);

ninexnine_unit ninexnine_unit_2926(
				.clk(clk),
				.rstn(rstn),
				.a0(P1221),
				.a1(P1231),
				.a2(P1241),
				.a3(P1321),
				.a4(P1331),
				.a5(P1341),
				.a6(P1421),
				.a7(P1431),
				.a8(P1441),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1122F)
);

ninexnine_unit ninexnine_unit_2927(
				.clk(clk),
				.rstn(rstn),
				.a0(P1222),
				.a1(P1232),
				.a2(P1242),
				.a3(P1322),
				.a4(P1332),
				.a5(P1342),
				.a6(P1422),
				.a7(P1432),
				.a8(P1442),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1222F)
);

assign C122F=c1022F+c1122F+c1222F;
assign A122F=(C122F>=0)?1:0;

assign P222F=A122F;

ninexnine_unit ninexnine_unit_2928(
				.clk(clk),
				.rstn(rstn),
				.a0(P1230),
				.a1(P1240),
				.a2(P1250),
				.a3(P1330),
				.a4(P1340),
				.a5(P1350),
				.a6(P1430),
				.a7(P1440),
				.a8(P1450),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1023F)
);

ninexnine_unit ninexnine_unit_2929(
				.clk(clk),
				.rstn(rstn),
				.a0(P1231),
				.a1(P1241),
				.a2(P1251),
				.a3(P1331),
				.a4(P1341),
				.a5(P1351),
				.a6(P1431),
				.a7(P1441),
				.a8(P1451),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1123F)
);

ninexnine_unit ninexnine_unit_2930(
				.clk(clk),
				.rstn(rstn),
				.a0(P1232),
				.a1(P1242),
				.a2(P1252),
				.a3(P1332),
				.a4(P1342),
				.a5(P1352),
				.a6(P1432),
				.a7(P1442),
				.a8(P1452),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1223F)
);

assign C123F=c1023F+c1123F+c1223F;
assign A123F=(C123F>=0)?1:0;

assign P223F=A123F;

ninexnine_unit ninexnine_unit_2931(
				.clk(clk),
				.rstn(rstn),
				.a0(P1240),
				.a1(P1250),
				.a2(P1260),
				.a3(P1340),
				.a4(P1350),
				.a5(P1360),
				.a6(P1440),
				.a7(P1450),
				.a8(P1460),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1024F)
);

ninexnine_unit ninexnine_unit_2932(
				.clk(clk),
				.rstn(rstn),
				.a0(P1241),
				.a1(P1251),
				.a2(P1261),
				.a3(P1341),
				.a4(P1351),
				.a5(P1361),
				.a6(P1441),
				.a7(P1451),
				.a8(P1461),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1124F)
);

ninexnine_unit ninexnine_unit_2933(
				.clk(clk),
				.rstn(rstn),
				.a0(P1242),
				.a1(P1252),
				.a2(P1262),
				.a3(P1342),
				.a4(P1352),
				.a5(P1362),
				.a6(P1442),
				.a7(P1452),
				.a8(P1462),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1224F)
);

assign C124F=c1024F+c1124F+c1224F;
assign A124F=(C124F>=0)?1:0;

assign P224F=A124F;

ninexnine_unit ninexnine_unit_2934(
				.clk(clk),
				.rstn(rstn),
				.a0(P1300),
				.a1(P1310),
				.a2(P1320),
				.a3(P1400),
				.a4(P1410),
				.a5(P1420),
				.a6(P1500),
				.a7(P1510),
				.a8(P1520),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1030F)
);

ninexnine_unit ninexnine_unit_2935(
				.clk(clk),
				.rstn(rstn),
				.a0(P1301),
				.a1(P1311),
				.a2(P1321),
				.a3(P1401),
				.a4(P1411),
				.a5(P1421),
				.a6(P1501),
				.a7(P1511),
				.a8(P1521),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1130F)
);

ninexnine_unit ninexnine_unit_2936(
				.clk(clk),
				.rstn(rstn),
				.a0(P1302),
				.a1(P1312),
				.a2(P1322),
				.a3(P1402),
				.a4(P1412),
				.a5(P1422),
				.a6(P1502),
				.a7(P1512),
				.a8(P1522),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1230F)
);

assign C130F=c1030F+c1130F+c1230F;
assign A130F=(C130F>=0)?1:0;

assign P230F=A130F;

ninexnine_unit ninexnine_unit_2937(
				.clk(clk),
				.rstn(rstn),
				.a0(P1310),
				.a1(P1320),
				.a2(P1330),
				.a3(P1410),
				.a4(P1420),
				.a5(P1430),
				.a6(P1510),
				.a7(P1520),
				.a8(P1530),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1031F)
);

ninexnine_unit ninexnine_unit_2938(
				.clk(clk),
				.rstn(rstn),
				.a0(P1311),
				.a1(P1321),
				.a2(P1331),
				.a3(P1411),
				.a4(P1421),
				.a5(P1431),
				.a6(P1511),
				.a7(P1521),
				.a8(P1531),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1131F)
);

ninexnine_unit ninexnine_unit_2939(
				.clk(clk),
				.rstn(rstn),
				.a0(P1312),
				.a1(P1322),
				.a2(P1332),
				.a3(P1412),
				.a4(P1422),
				.a5(P1432),
				.a6(P1512),
				.a7(P1522),
				.a8(P1532),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1231F)
);

assign C131F=c1031F+c1131F+c1231F;
assign A131F=(C131F>=0)?1:0;

assign P231F=A131F;

ninexnine_unit ninexnine_unit_2940(
				.clk(clk),
				.rstn(rstn),
				.a0(P1320),
				.a1(P1330),
				.a2(P1340),
				.a3(P1420),
				.a4(P1430),
				.a5(P1440),
				.a6(P1520),
				.a7(P1530),
				.a8(P1540),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1032F)
);

ninexnine_unit ninexnine_unit_2941(
				.clk(clk),
				.rstn(rstn),
				.a0(P1321),
				.a1(P1331),
				.a2(P1341),
				.a3(P1421),
				.a4(P1431),
				.a5(P1441),
				.a6(P1521),
				.a7(P1531),
				.a8(P1541),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1132F)
);

ninexnine_unit ninexnine_unit_2942(
				.clk(clk),
				.rstn(rstn),
				.a0(P1322),
				.a1(P1332),
				.a2(P1342),
				.a3(P1422),
				.a4(P1432),
				.a5(P1442),
				.a6(P1522),
				.a7(P1532),
				.a8(P1542),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1232F)
);

assign C132F=c1032F+c1132F+c1232F;
assign A132F=(C132F>=0)?1:0;

assign P232F=A132F;

ninexnine_unit ninexnine_unit_2943(
				.clk(clk),
				.rstn(rstn),
				.a0(P1330),
				.a1(P1340),
				.a2(P1350),
				.a3(P1430),
				.a4(P1440),
				.a5(P1450),
				.a6(P1530),
				.a7(P1540),
				.a8(P1550),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1033F)
);

ninexnine_unit ninexnine_unit_2944(
				.clk(clk),
				.rstn(rstn),
				.a0(P1331),
				.a1(P1341),
				.a2(P1351),
				.a3(P1431),
				.a4(P1441),
				.a5(P1451),
				.a6(P1531),
				.a7(P1541),
				.a8(P1551),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1133F)
);

ninexnine_unit ninexnine_unit_2945(
				.clk(clk),
				.rstn(rstn),
				.a0(P1332),
				.a1(P1342),
				.a2(P1352),
				.a3(P1432),
				.a4(P1442),
				.a5(P1452),
				.a6(P1532),
				.a7(P1542),
				.a8(P1552),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1233F)
);

assign C133F=c1033F+c1133F+c1233F;
assign A133F=(C133F>=0)?1:0;

assign P233F=A133F;

ninexnine_unit ninexnine_unit_2946(
				.clk(clk),
				.rstn(rstn),
				.a0(P1340),
				.a1(P1350),
				.a2(P1360),
				.a3(P1440),
				.a4(P1450),
				.a5(P1460),
				.a6(P1540),
				.a7(P1550),
				.a8(P1560),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1034F)
);

ninexnine_unit ninexnine_unit_2947(
				.clk(clk),
				.rstn(rstn),
				.a0(P1341),
				.a1(P1351),
				.a2(P1361),
				.a3(P1441),
				.a4(P1451),
				.a5(P1461),
				.a6(P1541),
				.a7(P1551),
				.a8(P1561),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1134F)
);

ninexnine_unit ninexnine_unit_2948(
				.clk(clk),
				.rstn(rstn),
				.a0(P1342),
				.a1(P1352),
				.a2(P1362),
				.a3(P1442),
				.a4(P1452),
				.a5(P1462),
				.a6(P1542),
				.a7(P1552),
				.a8(P1562),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1234F)
);

assign C134F=c1034F+c1134F+c1234F;
assign A134F=(C134F>=0)?1:0;

assign P234F=A134F;

ninexnine_unit ninexnine_unit_2949(
				.clk(clk),
				.rstn(rstn),
				.a0(P1400),
				.a1(P1410),
				.a2(P1420),
				.a3(P1500),
				.a4(P1510),
				.a5(P1520),
				.a6(P1600),
				.a7(P1610),
				.a8(P1620),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1040F)
);

ninexnine_unit ninexnine_unit_2950(
				.clk(clk),
				.rstn(rstn),
				.a0(P1401),
				.a1(P1411),
				.a2(P1421),
				.a3(P1501),
				.a4(P1511),
				.a5(P1521),
				.a6(P1601),
				.a7(P1611),
				.a8(P1621),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1140F)
);

ninexnine_unit ninexnine_unit_2951(
				.clk(clk),
				.rstn(rstn),
				.a0(P1402),
				.a1(P1412),
				.a2(P1422),
				.a3(P1502),
				.a4(P1512),
				.a5(P1522),
				.a6(P1602),
				.a7(P1612),
				.a8(P1622),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1240F)
);

assign C140F=c1040F+c1140F+c1240F;
assign A140F=(C140F>=0)?1:0;

assign P240F=A140F;

ninexnine_unit ninexnine_unit_2952(
				.clk(clk),
				.rstn(rstn),
				.a0(P1410),
				.a1(P1420),
				.a2(P1430),
				.a3(P1510),
				.a4(P1520),
				.a5(P1530),
				.a6(P1610),
				.a7(P1620),
				.a8(P1630),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1041F)
);

ninexnine_unit ninexnine_unit_2953(
				.clk(clk),
				.rstn(rstn),
				.a0(P1411),
				.a1(P1421),
				.a2(P1431),
				.a3(P1511),
				.a4(P1521),
				.a5(P1531),
				.a6(P1611),
				.a7(P1621),
				.a8(P1631),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1141F)
);

ninexnine_unit ninexnine_unit_2954(
				.clk(clk),
				.rstn(rstn),
				.a0(P1412),
				.a1(P1422),
				.a2(P1432),
				.a3(P1512),
				.a4(P1522),
				.a5(P1532),
				.a6(P1612),
				.a7(P1622),
				.a8(P1632),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1241F)
);

assign C141F=c1041F+c1141F+c1241F;
assign A141F=(C141F>=0)?1:0;

assign P241F=A141F;

ninexnine_unit ninexnine_unit_2955(
				.clk(clk),
				.rstn(rstn),
				.a0(P1420),
				.a1(P1430),
				.a2(P1440),
				.a3(P1520),
				.a4(P1530),
				.a5(P1540),
				.a6(P1620),
				.a7(P1630),
				.a8(P1640),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1042F)
);

ninexnine_unit ninexnine_unit_2956(
				.clk(clk),
				.rstn(rstn),
				.a0(P1421),
				.a1(P1431),
				.a2(P1441),
				.a3(P1521),
				.a4(P1531),
				.a5(P1541),
				.a6(P1621),
				.a7(P1631),
				.a8(P1641),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1142F)
);

ninexnine_unit ninexnine_unit_2957(
				.clk(clk),
				.rstn(rstn),
				.a0(P1422),
				.a1(P1432),
				.a2(P1442),
				.a3(P1522),
				.a4(P1532),
				.a5(P1542),
				.a6(P1622),
				.a7(P1632),
				.a8(P1642),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1242F)
);

assign C142F=c1042F+c1142F+c1242F;
assign A142F=(C142F>=0)?1:0;

assign P242F=A142F;

ninexnine_unit ninexnine_unit_2958(
				.clk(clk),
				.rstn(rstn),
				.a0(P1430),
				.a1(P1440),
				.a2(P1450),
				.a3(P1530),
				.a4(P1540),
				.a5(P1550),
				.a6(P1630),
				.a7(P1640),
				.a8(P1650),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1043F)
);

ninexnine_unit ninexnine_unit_2959(
				.clk(clk),
				.rstn(rstn),
				.a0(P1431),
				.a1(P1441),
				.a2(P1451),
				.a3(P1531),
				.a4(P1541),
				.a5(P1551),
				.a6(P1631),
				.a7(P1641),
				.a8(P1651),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1143F)
);

ninexnine_unit ninexnine_unit_2960(
				.clk(clk),
				.rstn(rstn),
				.a0(P1432),
				.a1(P1442),
				.a2(P1452),
				.a3(P1532),
				.a4(P1542),
				.a5(P1552),
				.a6(P1632),
				.a7(P1642),
				.a8(P1652),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1243F)
);

assign C143F=c1043F+c1143F+c1243F;
assign A143F=(C143F>=0)?1:0;

assign P243F=A143F;

ninexnine_unit ninexnine_unit_2961(
				.clk(clk),
				.rstn(rstn),
				.a0(P1440),
				.a1(P1450),
				.a2(P1460),
				.a3(P1540),
				.a4(P1550),
				.a5(P1560),
				.a6(P1640),
				.a7(P1650),
				.a8(P1660),
				.b0(W1F000),
				.b1(W1F010),
				.b2(W1F020),
				.b3(W1F100),
				.b4(W1F110),
				.b5(W1F120),
				.b6(W1F200),
				.b7(W1F210),
				.b8(W1F220),
				.c(c1044F)
);

ninexnine_unit ninexnine_unit_2962(
				.clk(clk),
				.rstn(rstn),
				.a0(P1441),
				.a1(P1451),
				.a2(P1461),
				.a3(P1541),
				.a4(P1551),
				.a5(P1561),
				.a6(P1641),
				.a7(P1651),
				.a8(P1661),
				.b0(W1F001),
				.b1(W1F011),
				.b2(W1F021),
				.b3(W1F101),
				.b4(W1F111),
				.b5(W1F121),
				.b6(W1F201),
				.b7(W1F211),
				.b8(W1F221),
				.c(c1144F)
);

ninexnine_unit ninexnine_unit_2963(
				.clk(clk),
				.rstn(rstn),
				.a0(P1442),
				.a1(P1452),
				.a2(P1462),
				.a3(P1542),
				.a4(P1552),
				.a5(P1562),
				.a6(P1642),
				.a7(P1652),
				.a8(P1662),
				.b0(W1F002),
				.b1(W1F012),
				.b2(W1F022),
				.b3(W1F102),
				.b4(W1F112),
				.b5(W1F122),
				.b6(W1F202),
				.b7(W1F212),
				.b8(W1F222),
				.c(c1244F)
);

assign C144F=c1044F+c1144F+c1244F;
assign A144F=(C144F>=0)?1:0;

assign P244F=A144F;

//layer2 done, begain next layer
wire P3000;
wire P3010;
wire P3020;
wire P3100;
wire P3110;
wire P3120;
wire P3200;
wire P3210;
wire P3220;
wire P3001;
wire P3011;
wire P3021;
wire P3101;
wire P3111;
wire P3121;
wire P3201;
wire P3211;
wire P3221;
wire P3002;
wire P3012;
wire P3022;
wire P3102;
wire P3112;
wire P3122;
wire P3202;
wire P3212;
wire P3222;
wire P3003;
wire P3013;
wire P3023;
wire P3103;
wire P3113;
wire P3123;
wire P3203;
wire P3213;
wire P3223;
wire P3004;
wire P3014;
wire P3024;
wire P3104;
wire P3114;
wire P3124;
wire P3204;
wire P3214;
wire P3224;
wire P3005;
wire P3015;
wire P3025;
wire P3105;
wire P3115;
wire P3125;
wire P3205;
wire P3215;
wire P3225;
wire P3006;
wire P3016;
wire P3026;
wire P3106;
wire P3116;
wire P3126;
wire P3206;
wire P3216;
wire P3226;
wire P3007;
wire P3017;
wire P3027;
wire P3107;
wire P3117;
wire P3127;
wire P3207;
wire P3217;
wire P3227;
wire P3008;
wire P3018;
wire P3028;
wire P3108;
wire P3118;
wire P3128;
wire P3208;
wire P3218;
wire P3228;
wire P3009;
wire P3019;
wire P3029;
wire P3109;
wire P3119;
wire P3129;
wire P3209;
wire P3219;
wire P3229;
wire P300A;
wire P301A;
wire P302A;
wire P310A;
wire P311A;
wire P312A;
wire P320A;
wire P321A;
wire P322A;
wire P300B;
wire P301B;
wire P302B;
wire P310B;
wire P311B;
wire P312B;
wire P320B;
wire P321B;
wire P322B;
wire P300C;
wire P301C;
wire P302C;
wire P310C;
wire P311C;
wire P312C;
wire P320C;
wire P321C;
wire P322C;
wire P300D;
wire P301D;
wire P302D;
wire P310D;
wire P311D;
wire P312D;
wire P320D;
wire P321D;
wire P322D;
wire P300E;
wire P301E;
wire P302E;
wire P310E;
wire P311E;
wire P312E;
wire P320E;
wire P321E;
wire P322E;
wire P300F;
wire P301F;
wire P302F;
wire P310F;
wire P311F;
wire P312F;
wire P320F;
wire P321F;
wire P322F;
wire P300G;
wire P301G;
wire P302G;
wire P310G;
wire P311G;
wire P312G;
wire P320G;
wire P321G;
wire P322G;
wire P300H;
wire P301H;
wire P302H;
wire P310H;
wire P311H;
wire P312H;
wire P320H;
wire P321H;
wire P322H;
wire P300I;
wire P301I;
wire P302I;
wire P310I;
wire P311I;
wire P312I;
wire P320I;
wire P321I;
wire P322I;
wire P300J;
wire P301J;
wire P302J;
wire P310J;
wire P311J;
wire P312J;
wire P320J;
wire P321J;
wire P322J;
wire P300K;
wire P301K;
wire P302K;
wire P310K;
wire P311K;
wire P312K;
wire P320K;
wire P321K;
wire P322K;
wire P300L;
wire P301L;
wire P302L;
wire P310L;
wire P311L;
wire P312L;
wire P320L;
wire P321L;
wire P322L;
wire P300M;
wire P301M;
wire P302M;
wire P310M;
wire P311M;
wire P312M;
wire P320M;
wire P321M;
wire P322M;
wire P300N;
wire P301N;
wire P302N;
wire P310N;
wire P311N;
wire P312N;
wire P320N;
wire P321N;
wire P322N;
wire P300O;
wire P301O;
wire P302O;
wire P310O;
wire P311O;
wire P312O;
wire P320O;
wire P321O;
wire P322O;
wire P300P;
wire P301P;
wire P302P;
wire P310P;
wire P311P;
wire P312P;
wire P320P;
wire P321P;
wire P322P;
wire P300Q;
wire P301Q;
wire P302Q;
wire P310Q;
wire P311Q;
wire P312Q;
wire P320Q;
wire P321Q;
wire P322Q;
wire P300R;
wire P301R;
wire P302R;
wire P310R;
wire P311R;
wire P312R;
wire P320R;
wire P321R;
wire P322R;
wire P300S;
wire P301S;
wire P302S;
wire P310S;
wire P311S;
wire P312S;
wire P320S;
wire P321S;
wire P322S;
wire P300T;
wire P301T;
wire P302T;
wire P310T;
wire P311T;
wire P312T;
wire P320T;
wire P321T;
wire P322T;
wire P300U;
wire P301U;
wire P302U;
wire P310U;
wire P311U;
wire P312U;
wire P320U;
wire P321U;
wire P322U;
wire P300V;
wire P301V;
wire P302V;
wire P310V;
wire P311V;
wire P312V;
wire P320V;
wire P321V;
wire P322V;
wire W20000,W20010,W20020,W20100,W20110,W20120,W20200,W20210,W20220;
wire W20001,W20011,W20021,W20101,W20111,W20121,W20201,W20211,W20221;
wire W20002,W20012,W20022,W20102,W20112,W20122,W20202,W20212,W20222;
wire W20003,W20013,W20023,W20103,W20113,W20123,W20203,W20213,W20223;
wire W20004,W20014,W20024,W20104,W20114,W20124,W20204,W20214,W20224;
wire W20005,W20015,W20025,W20105,W20115,W20125,W20205,W20215,W20225;
wire W20006,W20016,W20026,W20106,W20116,W20126,W20206,W20216,W20226;
wire W20007,W20017,W20027,W20107,W20117,W20127,W20207,W20217,W20227;
wire W20008,W20018,W20028,W20108,W20118,W20128,W20208,W20218,W20228;
wire W20009,W20019,W20029,W20109,W20119,W20129,W20209,W20219,W20229;
wire W2000A,W2001A,W2002A,W2010A,W2011A,W2012A,W2020A,W2021A,W2022A;
wire W2000B,W2001B,W2002B,W2010B,W2011B,W2012B,W2020B,W2021B,W2022B;
wire W2000C,W2001C,W2002C,W2010C,W2011C,W2012C,W2020C,W2021C,W2022C;
wire W2000D,W2001D,W2002D,W2010D,W2011D,W2012D,W2020D,W2021D,W2022D;
wire W2000E,W2001E,W2002E,W2010E,W2011E,W2012E,W2020E,W2021E,W2022E;
wire W2000F,W2001F,W2002F,W2010F,W2011F,W2012F,W2020F,W2021F,W2022F;
wire W21000,W21010,W21020,W21100,W21110,W21120,W21200,W21210,W21220;
wire W21001,W21011,W21021,W21101,W21111,W21121,W21201,W21211,W21221;
wire W21002,W21012,W21022,W21102,W21112,W21122,W21202,W21212,W21222;
wire W21003,W21013,W21023,W21103,W21113,W21123,W21203,W21213,W21223;
wire W21004,W21014,W21024,W21104,W21114,W21124,W21204,W21214,W21224;
wire W21005,W21015,W21025,W21105,W21115,W21125,W21205,W21215,W21225;
wire W21006,W21016,W21026,W21106,W21116,W21126,W21206,W21216,W21226;
wire W21007,W21017,W21027,W21107,W21117,W21127,W21207,W21217,W21227;
wire W21008,W21018,W21028,W21108,W21118,W21128,W21208,W21218,W21228;
wire W21009,W21019,W21029,W21109,W21119,W21129,W21209,W21219,W21229;
wire W2100A,W2101A,W2102A,W2110A,W2111A,W2112A,W2120A,W2121A,W2122A;
wire W2100B,W2101B,W2102B,W2110B,W2111B,W2112B,W2120B,W2121B,W2122B;
wire W2100C,W2101C,W2102C,W2110C,W2111C,W2112C,W2120C,W2121C,W2122C;
wire W2100D,W2101D,W2102D,W2110D,W2111D,W2112D,W2120D,W2121D,W2122D;
wire W2100E,W2101E,W2102E,W2110E,W2111E,W2112E,W2120E,W2121E,W2122E;
wire W2100F,W2101F,W2102F,W2110F,W2111F,W2112F,W2120F,W2121F,W2122F;
wire W22000,W22010,W22020,W22100,W22110,W22120,W22200,W22210,W22220;
wire W22001,W22011,W22021,W22101,W22111,W22121,W22201,W22211,W22221;
wire W22002,W22012,W22022,W22102,W22112,W22122,W22202,W22212,W22222;
wire W22003,W22013,W22023,W22103,W22113,W22123,W22203,W22213,W22223;
wire W22004,W22014,W22024,W22104,W22114,W22124,W22204,W22214,W22224;
wire W22005,W22015,W22025,W22105,W22115,W22125,W22205,W22215,W22225;
wire W22006,W22016,W22026,W22106,W22116,W22126,W22206,W22216,W22226;
wire W22007,W22017,W22027,W22107,W22117,W22127,W22207,W22217,W22227;
wire W22008,W22018,W22028,W22108,W22118,W22128,W22208,W22218,W22228;
wire W22009,W22019,W22029,W22109,W22119,W22129,W22209,W22219,W22229;
wire W2200A,W2201A,W2202A,W2210A,W2211A,W2212A,W2220A,W2221A,W2222A;
wire W2200B,W2201B,W2202B,W2210B,W2211B,W2212B,W2220B,W2221B,W2222B;
wire W2200C,W2201C,W2202C,W2210C,W2211C,W2212C,W2220C,W2221C,W2222C;
wire W2200D,W2201D,W2202D,W2210D,W2211D,W2212D,W2220D,W2221D,W2222D;
wire W2200E,W2201E,W2202E,W2210E,W2211E,W2212E,W2220E,W2221E,W2222E;
wire W2200F,W2201F,W2202F,W2210F,W2211F,W2212F,W2220F,W2221F,W2222F;
wire W23000,W23010,W23020,W23100,W23110,W23120,W23200,W23210,W23220;
wire W23001,W23011,W23021,W23101,W23111,W23121,W23201,W23211,W23221;
wire W23002,W23012,W23022,W23102,W23112,W23122,W23202,W23212,W23222;
wire W23003,W23013,W23023,W23103,W23113,W23123,W23203,W23213,W23223;
wire W23004,W23014,W23024,W23104,W23114,W23124,W23204,W23214,W23224;
wire W23005,W23015,W23025,W23105,W23115,W23125,W23205,W23215,W23225;
wire W23006,W23016,W23026,W23106,W23116,W23126,W23206,W23216,W23226;
wire W23007,W23017,W23027,W23107,W23117,W23127,W23207,W23217,W23227;
wire W23008,W23018,W23028,W23108,W23118,W23128,W23208,W23218,W23228;
wire W23009,W23019,W23029,W23109,W23119,W23129,W23209,W23219,W23229;
wire W2300A,W2301A,W2302A,W2310A,W2311A,W2312A,W2320A,W2321A,W2322A;
wire W2300B,W2301B,W2302B,W2310B,W2311B,W2312B,W2320B,W2321B,W2322B;
wire W2300C,W2301C,W2302C,W2310C,W2311C,W2312C,W2320C,W2321C,W2322C;
wire W2300D,W2301D,W2302D,W2310D,W2311D,W2312D,W2320D,W2321D,W2322D;
wire W2300E,W2301E,W2302E,W2310E,W2311E,W2312E,W2320E,W2321E,W2322E;
wire W2300F,W2301F,W2302F,W2310F,W2311F,W2312F,W2320F,W2321F,W2322F;
wire W24000,W24010,W24020,W24100,W24110,W24120,W24200,W24210,W24220;
wire W24001,W24011,W24021,W24101,W24111,W24121,W24201,W24211,W24221;
wire W24002,W24012,W24022,W24102,W24112,W24122,W24202,W24212,W24222;
wire W24003,W24013,W24023,W24103,W24113,W24123,W24203,W24213,W24223;
wire W24004,W24014,W24024,W24104,W24114,W24124,W24204,W24214,W24224;
wire W24005,W24015,W24025,W24105,W24115,W24125,W24205,W24215,W24225;
wire W24006,W24016,W24026,W24106,W24116,W24126,W24206,W24216,W24226;
wire W24007,W24017,W24027,W24107,W24117,W24127,W24207,W24217,W24227;
wire W24008,W24018,W24028,W24108,W24118,W24128,W24208,W24218,W24228;
wire W24009,W24019,W24029,W24109,W24119,W24129,W24209,W24219,W24229;
wire W2400A,W2401A,W2402A,W2410A,W2411A,W2412A,W2420A,W2421A,W2422A;
wire W2400B,W2401B,W2402B,W2410B,W2411B,W2412B,W2420B,W2421B,W2422B;
wire W2400C,W2401C,W2402C,W2410C,W2411C,W2412C,W2420C,W2421C,W2422C;
wire W2400D,W2401D,W2402D,W2410D,W2411D,W2412D,W2420D,W2421D,W2422D;
wire W2400E,W2401E,W2402E,W2410E,W2411E,W2412E,W2420E,W2421E,W2422E;
wire W2400F,W2401F,W2402F,W2410F,W2411F,W2412F,W2420F,W2421F,W2422F;
wire W25000,W25010,W25020,W25100,W25110,W25120,W25200,W25210,W25220;
wire W25001,W25011,W25021,W25101,W25111,W25121,W25201,W25211,W25221;
wire W25002,W25012,W25022,W25102,W25112,W25122,W25202,W25212,W25222;
wire W25003,W25013,W25023,W25103,W25113,W25123,W25203,W25213,W25223;
wire W25004,W25014,W25024,W25104,W25114,W25124,W25204,W25214,W25224;
wire W25005,W25015,W25025,W25105,W25115,W25125,W25205,W25215,W25225;
wire W25006,W25016,W25026,W25106,W25116,W25126,W25206,W25216,W25226;
wire W25007,W25017,W25027,W25107,W25117,W25127,W25207,W25217,W25227;
wire W25008,W25018,W25028,W25108,W25118,W25128,W25208,W25218,W25228;
wire W25009,W25019,W25029,W25109,W25119,W25129,W25209,W25219,W25229;
wire W2500A,W2501A,W2502A,W2510A,W2511A,W2512A,W2520A,W2521A,W2522A;
wire W2500B,W2501B,W2502B,W2510B,W2511B,W2512B,W2520B,W2521B,W2522B;
wire W2500C,W2501C,W2502C,W2510C,W2511C,W2512C,W2520C,W2521C,W2522C;
wire W2500D,W2501D,W2502D,W2510D,W2511D,W2512D,W2520D,W2521D,W2522D;
wire W2500E,W2501E,W2502E,W2510E,W2511E,W2512E,W2520E,W2521E,W2522E;
wire W2500F,W2501F,W2502F,W2510F,W2511F,W2512F,W2520F,W2521F,W2522F;
wire W26000,W26010,W26020,W26100,W26110,W26120,W26200,W26210,W26220;
wire W26001,W26011,W26021,W26101,W26111,W26121,W26201,W26211,W26221;
wire W26002,W26012,W26022,W26102,W26112,W26122,W26202,W26212,W26222;
wire W26003,W26013,W26023,W26103,W26113,W26123,W26203,W26213,W26223;
wire W26004,W26014,W26024,W26104,W26114,W26124,W26204,W26214,W26224;
wire W26005,W26015,W26025,W26105,W26115,W26125,W26205,W26215,W26225;
wire W26006,W26016,W26026,W26106,W26116,W26126,W26206,W26216,W26226;
wire W26007,W26017,W26027,W26107,W26117,W26127,W26207,W26217,W26227;
wire W26008,W26018,W26028,W26108,W26118,W26128,W26208,W26218,W26228;
wire W26009,W26019,W26029,W26109,W26119,W26129,W26209,W26219,W26229;
wire W2600A,W2601A,W2602A,W2610A,W2611A,W2612A,W2620A,W2621A,W2622A;
wire W2600B,W2601B,W2602B,W2610B,W2611B,W2612B,W2620B,W2621B,W2622B;
wire W2600C,W2601C,W2602C,W2610C,W2611C,W2612C,W2620C,W2621C,W2622C;
wire W2600D,W2601D,W2602D,W2610D,W2611D,W2612D,W2620D,W2621D,W2622D;
wire W2600E,W2601E,W2602E,W2610E,W2611E,W2612E,W2620E,W2621E,W2622E;
wire W2600F,W2601F,W2602F,W2610F,W2611F,W2612F,W2620F,W2621F,W2622F;
wire W27000,W27010,W27020,W27100,W27110,W27120,W27200,W27210,W27220;
wire W27001,W27011,W27021,W27101,W27111,W27121,W27201,W27211,W27221;
wire W27002,W27012,W27022,W27102,W27112,W27122,W27202,W27212,W27222;
wire W27003,W27013,W27023,W27103,W27113,W27123,W27203,W27213,W27223;
wire W27004,W27014,W27024,W27104,W27114,W27124,W27204,W27214,W27224;
wire W27005,W27015,W27025,W27105,W27115,W27125,W27205,W27215,W27225;
wire W27006,W27016,W27026,W27106,W27116,W27126,W27206,W27216,W27226;
wire W27007,W27017,W27027,W27107,W27117,W27127,W27207,W27217,W27227;
wire W27008,W27018,W27028,W27108,W27118,W27128,W27208,W27218,W27228;
wire W27009,W27019,W27029,W27109,W27119,W27129,W27209,W27219,W27229;
wire W2700A,W2701A,W2702A,W2710A,W2711A,W2712A,W2720A,W2721A,W2722A;
wire W2700B,W2701B,W2702B,W2710B,W2711B,W2712B,W2720B,W2721B,W2722B;
wire W2700C,W2701C,W2702C,W2710C,W2711C,W2712C,W2720C,W2721C,W2722C;
wire W2700D,W2701D,W2702D,W2710D,W2711D,W2712D,W2720D,W2721D,W2722D;
wire W2700E,W2701E,W2702E,W2710E,W2711E,W2712E,W2720E,W2721E,W2722E;
wire W2700F,W2701F,W2702F,W2710F,W2711F,W2712F,W2720F,W2721F,W2722F;
wire W28000,W28010,W28020,W28100,W28110,W28120,W28200,W28210,W28220;
wire W28001,W28011,W28021,W28101,W28111,W28121,W28201,W28211,W28221;
wire W28002,W28012,W28022,W28102,W28112,W28122,W28202,W28212,W28222;
wire W28003,W28013,W28023,W28103,W28113,W28123,W28203,W28213,W28223;
wire W28004,W28014,W28024,W28104,W28114,W28124,W28204,W28214,W28224;
wire W28005,W28015,W28025,W28105,W28115,W28125,W28205,W28215,W28225;
wire W28006,W28016,W28026,W28106,W28116,W28126,W28206,W28216,W28226;
wire W28007,W28017,W28027,W28107,W28117,W28127,W28207,W28217,W28227;
wire W28008,W28018,W28028,W28108,W28118,W28128,W28208,W28218,W28228;
wire W28009,W28019,W28029,W28109,W28119,W28129,W28209,W28219,W28229;
wire W2800A,W2801A,W2802A,W2810A,W2811A,W2812A,W2820A,W2821A,W2822A;
wire W2800B,W2801B,W2802B,W2810B,W2811B,W2812B,W2820B,W2821B,W2822B;
wire W2800C,W2801C,W2802C,W2810C,W2811C,W2812C,W2820C,W2821C,W2822C;
wire W2800D,W2801D,W2802D,W2810D,W2811D,W2812D,W2820D,W2821D,W2822D;
wire W2800E,W2801E,W2802E,W2810E,W2811E,W2812E,W2820E,W2821E,W2822E;
wire W2800F,W2801F,W2802F,W2810F,W2811F,W2812F,W2820F,W2821F,W2822F;
wire W29000,W29010,W29020,W29100,W29110,W29120,W29200,W29210,W29220;
wire W29001,W29011,W29021,W29101,W29111,W29121,W29201,W29211,W29221;
wire W29002,W29012,W29022,W29102,W29112,W29122,W29202,W29212,W29222;
wire W29003,W29013,W29023,W29103,W29113,W29123,W29203,W29213,W29223;
wire W29004,W29014,W29024,W29104,W29114,W29124,W29204,W29214,W29224;
wire W29005,W29015,W29025,W29105,W29115,W29125,W29205,W29215,W29225;
wire W29006,W29016,W29026,W29106,W29116,W29126,W29206,W29216,W29226;
wire W29007,W29017,W29027,W29107,W29117,W29127,W29207,W29217,W29227;
wire W29008,W29018,W29028,W29108,W29118,W29128,W29208,W29218,W29228;
wire W29009,W29019,W29029,W29109,W29119,W29129,W29209,W29219,W29229;
wire W2900A,W2901A,W2902A,W2910A,W2911A,W2912A,W2920A,W2921A,W2922A;
wire W2900B,W2901B,W2902B,W2910B,W2911B,W2912B,W2920B,W2921B,W2922B;
wire W2900C,W2901C,W2902C,W2910C,W2911C,W2912C,W2920C,W2921C,W2922C;
wire W2900D,W2901D,W2902D,W2910D,W2911D,W2912D,W2920D,W2921D,W2922D;
wire W2900E,W2901E,W2902E,W2910E,W2911E,W2912E,W2920E,W2921E,W2922E;
wire W2900F,W2901F,W2902F,W2910F,W2911F,W2912F,W2920F,W2921F,W2922F;
wire W2A000,W2A010,W2A020,W2A100,W2A110,W2A120,W2A200,W2A210,W2A220;
wire W2A001,W2A011,W2A021,W2A101,W2A111,W2A121,W2A201,W2A211,W2A221;
wire W2A002,W2A012,W2A022,W2A102,W2A112,W2A122,W2A202,W2A212,W2A222;
wire W2A003,W2A013,W2A023,W2A103,W2A113,W2A123,W2A203,W2A213,W2A223;
wire W2A004,W2A014,W2A024,W2A104,W2A114,W2A124,W2A204,W2A214,W2A224;
wire W2A005,W2A015,W2A025,W2A105,W2A115,W2A125,W2A205,W2A215,W2A225;
wire W2A006,W2A016,W2A026,W2A106,W2A116,W2A126,W2A206,W2A216,W2A226;
wire W2A007,W2A017,W2A027,W2A107,W2A117,W2A127,W2A207,W2A217,W2A227;
wire W2A008,W2A018,W2A028,W2A108,W2A118,W2A128,W2A208,W2A218,W2A228;
wire W2A009,W2A019,W2A029,W2A109,W2A119,W2A129,W2A209,W2A219,W2A229;
wire W2A00A,W2A01A,W2A02A,W2A10A,W2A11A,W2A12A,W2A20A,W2A21A,W2A22A;
wire W2A00B,W2A01B,W2A02B,W2A10B,W2A11B,W2A12B,W2A20B,W2A21B,W2A22B;
wire W2A00C,W2A01C,W2A02C,W2A10C,W2A11C,W2A12C,W2A20C,W2A21C,W2A22C;
wire W2A00D,W2A01D,W2A02D,W2A10D,W2A11D,W2A12D,W2A20D,W2A21D,W2A22D;
wire W2A00E,W2A01E,W2A02E,W2A10E,W2A11E,W2A12E,W2A20E,W2A21E,W2A22E;
wire W2A00F,W2A01F,W2A02F,W2A10F,W2A11F,W2A12F,W2A20F,W2A21F,W2A22F;
wire W2B000,W2B010,W2B020,W2B100,W2B110,W2B120,W2B200,W2B210,W2B220;
wire W2B001,W2B011,W2B021,W2B101,W2B111,W2B121,W2B201,W2B211,W2B221;
wire W2B002,W2B012,W2B022,W2B102,W2B112,W2B122,W2B202,W2B212,W2B222;
wire W2B003,W2B013,W2B023,W2B103,W2B113,W2B123,W2B203,W2B213,W2B223;
wire W2B004,W2B014,W2B024,W2B104,W2B114,W2B124,W2B204,W2B214,W2B224;
wire W2B005,W2B015,W2B025,W2B105,W2B115,W2B125,W2B205,W2B215,W2B225;
wire W2B006,W2B016,W2B026,W2B106,W2B116,W2B126,W2B206,W2B216,W2B226;
wire W2B007,W2B017,W2B027,W2B107,W2B117,W2B127,W2B207,W2B217,W2B227;
wire W2B008,W2B018,W2B028,W2B108,W2B118,W2B128,W2B208,W2B218,W2B228;
wire W2B009,W2B019,W2B029,W2B109,W2B119,W2B129,W2B209,W2B219,W2B229;
wire W2B00A,W2B01A,W2B02A,W2B10A,W2B11A,W2B12A,W2B20A,W2B21A,W2B22A;
wire W2B00B,W2B01B,W2B02B,W2B10B,W2B11B,W2B12B,W2B20B,W2B21B,W2B22B;
wire W2B00C,W2B01C,W2B02C,W2B10C,W2B11C,W2B12C,W2B20C,W2B21C,W2B22C;
wire W2B00D,W2B01D,W2B02D,W2B10D,W2B11D,W2B12D,W2B20D,W2B21D,W2B22D;
wire W2B00E,W2B01E,W2B02E,W2B10E,W2B11E,W2B12E,W2B20E,W2B21E,W2B22E;
wire W2B00F,W2B01F,W2B02F,W2B10F,W2B11F,W2B12F,W2B20F,W2B21F,W2B22F;
wire W2C000,W2C010,W2C020,W2C100,W2C110,W2C120,W2C200,W2C210,W2C220;
wire W2C001,W2C011,W2C021,W2C101,W2C111,W2C121,W2C201,W2C211,W2C221;
wire W2C002,W2C012,W2C022,W2C102,W2C112,W2C122,W2C202,W2C212,W2C222;
wire W2C003,W2C013,W2C023,W2C103,W2C113,W2C123,W2C203,W2C213,W2C223;
wire W2C004,W2C014,W2C024,W2C104,W2C114,W2C124,W2C204,W2C214,W2C224;
wire W2C005,W2C015,W2C025,W2C105,W2C115,W2C125,W2C205,W2C215,W2C225;
wire W2C006,W2C016,W2C026,W2C106,W2C116,W2C126,W2C206,W2C216,W2C226;
wire W2C007,W2C017,W2C027,W2C107,W2C117,W2C127,W2C207,W2C217,W2C227;
wire W2C008,W2C018,W2C028,W2C108,W2C118,W2C128,W2C208,W2C218,W2C228;
wire W2C009,W2C019,W2C029,W2C109,W2C119,W2C129,W2C209,W2C219,W2C229;
wire W2C00A,W2C01A,W2C02A,W2C10A,W2C11A,W2C12A,W2C20A,W2C21A,W2C22A;
wire W2C00B,W2C01B,W2C02B,W2C10B,W2C11B,W2C12B,W2C20B,W2C21B,W2C22B;
wire W2C00C,W2C01C,W2C02C,W2C10C,W2C11C,W2C12C,W2C20C,W2C21C,W2C22C;
wire W2C00D,W2C01D,W2C02D,W2C10D,W2C11D,W2C12D,W2C20D,W2C21D,W2C22D;
wire W2C00E,W2C01E,W2C02E,W2C10E,W2C11E,W2C12E,W2C20E,W2C21E,W2C22E;
wire W2C00F,W2C01F,W2C02F,W2C10F,W2C11F,W2C12F,W2C20F,W2C21F,W2C22F;
wire W2D000,W2D010,W2D020,W2D100,W2D110,W2D120,W2D200,W2D210,W2D220;
wire W2D001,W2D011,W2D021,W2D101,W2D111,W2D121,W2D201,W2D211,W2D221;
wire W2D002,W2D012,W2D022,W2D102,W2D112,W2D122,W2D202,W2D212,W2D222;
wire W2D003,W2D013,W2D023,W2D103,W2D113,W2D123,W2D203,W2D213,W2D223;
wire W2D004,W2D014,W2D024,W2D104,W2D114,W2D124,W2D204,W2D214,W2D224;
wire W2D005,W2D015,W2D025,W2D105,W2D115,W2D125,W2D205,W2D215,W2D225;
wire W2D006,W2D016,W2D026,W2D106,W2D116,W2D126,W2D206,W2D216,W2D226;
wire W2D007,W2D017,W2D027,W2D107,W2D117,W2D127,W2D207,W2D217,W2D227;
wire W2D008,W2D018,W2D028,W2D108,W2D118,W2D128,W2D208,W2D218,W2D228;
wire W2D009,W2D019,W2D029,W2D109,W2D119,W2D129,W2D209,W2D219,W2D229;
wire W2D00A,W2D01A,W2D02A,W2D10A,W2D11A,W2D12A,W2D20A,W2D21A,W2D22A;
wire W2D00B,W2D01B,W2D02B,W2D10B,W2D11B,W2D12B,W2D20B,W2D21B,W2D22B;
wire W2D00C,W2D01C,W2D02C,W2D10C,W2D11C,W2D12C,W2D20C,W2D21C,W2D22C;
wire W2D00D,W2D01D,W2D02D,W2D10D,W2D11D,W2D12D,W2D20D,W2D21D,W2D22D;
wire W2D00E,W2D01E,W2D02E,W2D10E,W2D11E,W2D12E,W2D20E,W2D21E,W2D22E;
wire W2D00F,W2D01F,W2D02F,W2D10F,W2D11F,W2D12F,W2D20F,W2D21F,W2D22F;
wire W2E000,W2E010,W2E020,W2E100,W2E110,W2E120,W2E200,W2E210,W2E220;
wire W2E001,W2E011,W2E021,W2E101,W2E111,W2E121,W2E201,W2E211,W2E221;
wire W2E002,W2E012,W2E022,W2E102,W2E112,W2E122,W2E202,W2E212,W2E222;
wire W2E003,W2E013,W2E023,W2E103,W2E113,W2E123,W2E203,W2E213,W2E223;
wire W2E004,W2E014,W2E024,W2E104,W2E114,W2E124,W2E204,W2E214,W2E224;
wire W2E005,W2E015,W2E025,W2E105,W2E115,W2E125,W2E205,W2E215,W2E225;
wire W2E006,W2E016,W2E026,W2E106,W2E116,W2E126,W2E206,W2E216,W2E226;
wire W2E007,W2E017,W2E027,W2E107,W2E117,W2E127,W2E207,W2E217,W2E227;
wire W2E008,W2E018,W2E028,W2E108,W2E118,W2E128,W2E208,W2E218,W2E228;
wire W2E009,W2E019,W2E029,W2E109,W2E119,W2E129,W2E209,W2E219,W2E229;
wire W2E00A,W2E01A,W2E02A,W2E10A,W2E11A,W2E12A,W2E20A,W2E21A,W2E22A;
wire W2E00B,W2E01B,W2E02B,W2E10B,W2E11B,W2E12B,W2E20B,W2E21B,W2E22B;
wire W2E00C,W2E01C,W2E02C,W2E10C,W2E11C,W2E12C,W2E20C,W2E21C,W2E22C;
wire W2E00D,W2E01D,W2E02D,W2E10D,W2E11D,W2E12D,W2E20D,W2E21D,W2E22D;
wire W2E00E,W2E01E,W2E02E,W2E10E,W2E11E,W2E12E,W2E20E,W2E21E,W2E22E;
wire W2E00F,W2E01F,W2E02F,W2E10F,W2E11F,W2E12F,W2E20F,W2E21F,W2E22F;
wire W2F000,W2F010,W2F020,W2F100,W2F110,W2F120,W2F200,W2F210,W2F220;
wire W2F001,W2F011,W2F021,W2F101,W2F111,W2F121,W2F201,W2F211,W2F221;
wire W2F002,W2F012,W2F022,W2F102,W2F112,W2F122,W2F202,W2F212,W2F222;
wire W2F003,W2F013,W2F023,W2F103,W2F113,W2F123,W2F203,W2F213,W2F223;
wire W2F004,W2F014,W2F024,W2F104,W2F114,W2F124,W2F204,W2F214,W2F224;
wire W2F005,W2F015,W2F025,W2F105,W2F115,W2F125,W2F205,W2F215,W2F225;
wire W2F006,W2F016,W2F026,W2F106,W2F116,W2F126,W2F206,W2F216,W2F226;
wire W2F007,W2F017,W2F027,W2F107,W2F117,W2F127,W2F207,W2F217,W2F227;
wire W2F008,W2F018,W2F028,W2F108,W2F118,W2F128,W2F208,W2F218,W2F228;
wire W2F009,W2F019,W2F029,W2F109,W2F119,W2F129,W2F209,W2F219,W2F229;
wire W2F00A,W2F01A,W2F02A,W2F10A,W2F11A,W2F12A,W2F20A,W2F21A,W2F22A;
wire W2F00B,W2F01B,W2F02B,W2F10B,W2F11B,W2F12B,W2F20B,W2F21B,W2F22B;
wire W2F00C,W2F01C,W2F02C,W2F10C,W2F11C,W2F12C,W2F20C,W2F21C,W2F22C;
wire W2F00D,W2F01D,W2F02D,W2F10D,W2F11D,W2F12D,W2F20D,W2F21D,W2F22D;
wire W2F00E,W2F01E,W2F02E,W2F10E,W2F11E,W2F12E,W2F20E,W2F21E,W2F22E;
wire W2F00F,W2F01F,W2F02F,W2F10F,W2F11F,W2F12F,W2F20F,W2F21F,W2F22F;
wire W2G000,W2G010,W2G020,W2G100,W2G110,W2G120,W2G200,W2G210,W2G220;
wire W2G001,W2G011,W2G021,W2G101,W2G111,W2G121,W2G201,W2G211,W2G221;
wire W2G002,W2G012,W2G022,W2G102,W2G112,W2G122,W2G202,W2G212,W2G222;
wire W2G003,W2G013,W2G023,W2G103,W2G113,W2G123,W2G203,W2G213,W2G223;
wire W2G004,W2G014,W2G024,W2G104,W2G114,W2G124,W2G204,W2G214,W2G224;
wire W2G005,W2G015,W2G025,W2G105,W2G115,W2G125,W2G205,W2G215,W2G225;
wire W2G006,W2G016,W2G026,W2G106,W2G116,W2G126,W2G206,W2G216,W2G226;
wire W2G007,W2G017,W2G027,W2G107,W2G117,W2G127,W2G207,W2G217,W2G227;
wire W2G008,W2G018,W2G028,W2G108,W2G118,W2G128,W2G208,W2G218,W2G228;
wire W2G009,W2G019,W2G029,W2G109,W2G119,W2G129,W2G209,W2G219,W2G229;
wire W2G00A,W2G01A,W2G02A,W2G10A,W2G11A,W2G12A,W2G20A,W2G21A,W2G22A;
wire W2G00B,W2G01B,W2G02B,W2G10B,W2G11B,W2G12B,W2G20B,W2G21B,W2G22B;
wire W2G00C,W2G01C,W2G02C,W2G10C,W2G11C,W2G12C,W2G20C,W2G21C,W2G22C;
wire W2G00D,W2G01D,W2G02D,W2G10D,W2G11D,W2G12D,W2G20D,W2G21D,W2G22D;
wire W2G00E,W2G01E,W2G02E,W2G10E,W2G11E,W2G12E,W2G20E,W2G21E,W2G22E;
wire W2G00F,W2G01F,W2G02F,W2G10F,W2G11F,W2G12F,W2G20F,W2G21F,W2G22F;
wire W2H000,W2H010,W2H020,W2H100,W2H110,W2H120,W2H200,W2H210,W2H220;
wire W2H001,W2H011,W2H021,W2H101,W2H111,W2H121,W2H201,W2H211,W2H221;
wire W2H002,W2H012,W2H022,W2H102,W2H112,W2H122,W2H202,W2H212,W2H222;
wire W2H003,W2H013,W2H023,W2H103,W2H113,W2H123,W2H203,W2H213,W2H223;
wire W2H004,W2H014,W2H024,W2H104,W2H114,W2H124,W2H204,W2H214,W2H224;
wire W2H005,W2H015,W2H025,W2H105,W2H115,W2H125,W2H205,W2H215,W2H225;
wire W2H006,W2H016,W2H026,W2H106,W2H116,W2H126,W2H206,W2H216,W2H226;
wire W2H007,W2H017,W2H027,W2H107,W2H117,W2H127,W2H207,W2H217,W2H227;
wire W2H008,W2H018,W2H028,W2H108,W2H118,W2H128,W2H208,W2H218,W2H228;
wire W2H009,W2H019,W2H029,W2H109,W2H119,W2H129,W2H209,W2H219,W2H229;
wire W2H00A,W2H01A,W2H02A,W2H10A,W2H11A,W2H12A,W2H20A,W2H21A,W2H22A;
wire W2H00B,W2H01B,W2H02B,W2H10B,W2H11B,W2H12B,W2H20B,W2H21B,W2H22B;
wire W2H00C,W2H01C,W2H02C,W2H10C,W2H11C,W2H12C,W2H20C,W2H21C,W2H22C;
wire W2H00D,W2H01D,W2H02D,W2H10D,W2H11D,W2H12D,W2H20D,W2H21D,W2H22D;
wire W2H00E,W2H01E,W2H02E,W2H10E,W2H11E,W2H12E,W2H20E,W2H21E,W2H22E;
wire W2H00F,W2H01F,W2H02F,W2H10F,W2H11F,W2H12F,W2H20F,W2H21F,W2H22F;
wire W2I000,W2I010,W2I020,W2I100,W2I110,W2I120,W2I200,W2I210,W2I220;
wire W2I001,W2I011,W2I021,W2I101,W2I111,W2I121,W2I201,W2I211,W2I221;
wire W2I002,W2I012,W2I022,W2I102,W2I112,W2I122,W2I202,W2I212,W2I222;
wire W2I003,W2I013,W2I023,W2I103,W2I113,W2I123,W2I203,W2I213,W2I223;
wire W2I004,W2I014,W2I024,W2I104,W2I114,W2I124,W2I204,W2I214,W2I224;
wire W2I005,W2I015,W2I025,W2I105,W2I115,W2I125,W2I205,W2I215,W2I225;
wire W2I006,W2I016,W2I026,W2I106,W2I116,W2I126,W2I206,W2I216,W2I226;
wire W2I007,W2I017,W2I027,W2I107,W2I117,W2I127,W2I207,W2I217,W2I227;
wire W2I008,W2I018,W2I028,W2I108,W2I118,W2I128,W2I208,W2I218,W2I228;
wire W2I009,W2I019,W2I029,W2I109,W2I119,W2I129,W2I209,W2I219,W2I229;
wire W2I00A,W2I01A,W2I02A,W2I10A,W2I11A,W2I12A,W2I20A,W2I21A,W2I22A;
wire W2I00B,W2I01B,W2I02B,W2I10B,W2I11B,W2I12B,W2I20B,W2I21B,W2I22B;
wire W2I00C,W2I01C,W2I02C,W2I10C,W2I11C,W2I12C,W2I20C,W2I21C,W2I22C;
wire W2I00D,W2I01D,W2I02D,W2I10D,W2I11D,W2I12D,W2I20D,W2I21D,W2I22D;
wire W2I00E,W2I01E,W2I02E,W2I10E,W2I11E,W2I12E,W2I20E,W2I21E,W2I22E;
wire W2I00F,W2I01F,W2I02F,W2I10F,W2I11F,W2I12F,W2I20F,W2I21F,W2I22F;
wire W2J000,W2J010,W2J020,W2J100,W2J110,W2J120,W2J200,W2J210,W2J220;
wire W2J001,W2J011,W2J021,W2J101,W2J111,W2J121,W2J201,W2J211,W2J221;
wire W2J002,W2J012,W2J022,W2J102,W2J112,W2J122,W2J202,W2J212,W2J222;
wire W2J003,W2J013,W2J023,W2J103,W2J113,W2J123,W2J203,W2J213,W2J223;
wire W2J004,W2J014,W2J024,W2J104,W2J114,W2J124,W2J204,W2J214,W2J224;
wire W2J005,W2J015,W2J025,W2J105,W2J115,W2J125,W2J205,W2J215,W2J225;
wire W2J006,W2J016,W2J026,W2J106,W2J116,W2J126,W2J206,W2J216,W2J226;
wire W2J007,W2J017,W2J027,W2J107,W2J117,W2J127,W2J207,W2J217,W2J227;
wire W2J008,W2J018,W2J028,W2J108,W2J118,W2J128,W2J208,W2J218,W2J228;
wire W2J009,W2J019,W2J029,W2J109,W2J119,W2J129,W2J209,W2J219,W2J229;
wire W2J00A,W2J01A,W2J02A,W2J10A,W2J11A,W2J12A,W2J20A,W2J21A,W2J22A;
wire W2J00B,W2J01B,W2J02B,W2J10B,W2J11B,W2J12B,W2J20B,W2J21B,W2J22B;
wire W2J00C,W2J01C,W2J02C,W2J10C,W2J11C,W2J12C,W2J20C,W2J21C,W2J22C;
wire W2J00D,W2J01D,W2J02D,W2J10D,W2J11D,W2J12D,W2J20D,W2J21D,W2J22D;
wire W2J00E,W2J01E,W2J02E,W2J10E,W2J11E,W2J12E,W2J20E,W2J21E,W2J22E;
wire W2J00F,W2J01F,W2J02F,W2J10F,W2J11F,W2J12F,W2J20F,W2J21F,W2J22F;
wire W2K000,W2K010,W2K020,W2K100,W2K110,W2K120,W2K200,W2K210,W2K220;
wire W2K001,W2K011,W2K021,W2K101,W2K111,W2K121,W2K201,W2K211,W2K221;
wire W2K002,W2K012,W2K022,W2K102,W2K112,W2K122,W2K202,W2K212,W2K222;
wire W2K003,W2K013,W2K023,W2K103,W2K113,W2K123,W2K203,W2K213,W2K223;
wire W2K004,W2K014,W2K024,W2K104,W2K114,W2K124,W2K204,W2K214,W2K224;
wire W2K005,W2K015,W2K025,W2K105,W2K115,W2K125,W2K205,W2K215,W2K225;
wire W2K006,W2K016,W2K026,W2K106,W2K116,W2K126,W2K206,W2K216,W2K226;
wire W2K007,W2K017,W2K027,W2K107,W2K117,W2K127,W2K207,W2K217,W2K227;
wire W2K008,W2K018,W2K028,W2K108,W2K118,W2K128,W2K208,W2K218,W2K228;
wire W2K009,W2K019,W2K029,W2K109,W2K119,W2K129,W2K209,W2K219,W2K229;
wire W2K00A,W2K01A,W2K02A,W2K10A,W2K11A,W2K12A,W2K20A,W2K21A,W2K22A;
wire W2K00B,W2K01B,W2K02B,W2K10B,W2K11B,W2K12B,W2K20B,W2K21B,W2K22B;
wire W2K00C,W2K01C,W2K02C,W2K10C,W2K11C,W2K12C,W2K20C,W2K21C,W2K22C;
wire W2K00D,W2K01D,W2K02D,W2K10D,W2K11D,W2K12D,W2K20D,W2K21D,W2K22D;
wire W2K00E,W2K01E,W2K02E,W2K10E,W2K11E,W2K12E,W2K20E,W2K21E,W2K22E;
wire W2K00F,W2K01F,W2K02F,W2K10F,W2K11F,W2K12F,W2K20F,W2K21F,W2K22F;
wire W2L000,W2L010,W2L020,W2L100,W2L110,W2L120,W2L200,W2L210,W2L220;
wire W2L001,W2L011,W2L021,W2L101,W2L111,W2L121,W2L201,W2L211,W2L221;
wire W2L002,W2L012,W2L022,W2L102,W2L112,W2L122,W2L202,W2L212,W2L222;
wire W2L003,W2L013,W2L023,W2L103,W2L113,W2L123,W2L203,W2L213,W2L223;
wire W2L004,W2L014,W2L024,W2L104,W2L114,W2L124,W2L204,W2L214,W2L224;
wire W2L005,W2L015,W2L025,W2L105,W2L115,W2L125,W2L205,W2L215,W2L225;
wire W2L006,W2L016,W2L026,W2L106,W2L116,W2L126,W2L206,W2L216,W2L226;
wire W2L007,W2L017,W2L027,W2L107,W2L117,W2L127,W2L207,W2L217,W2L227;
wire W2L008,W2L018,W2L028,W2L108,W2L118,W2L128,W2L208,W2L218,W2L228;
wire W2L009,W2L019,W2L029,W2L109,W2L119,W2L129,W2L209,W2L219,W2L229;
wire W2L00A,W2L01A,W2L02A,W2L10A,W2L11A,W2L12A,W2L20A,W2L21A,W2L22A;
wire W2L00B,W2L01B,W2L02B,W2L10B,W2L11B,W2L12B,W2L20B,W2L21B,W2L22B;
wire W2L00C,W2L01C,W2L02C,W2L10C,W2L11C,W2L12C,W2L20C,W2L21C,W2L22C;
wire W2L00D,W2L01D,W2L02D,W2L10D,W2L11D,W2L12D,W2L20D,W2L21D,W2L22D;
wire W2L00E,W2L01E,W2L02E,W2L10E,W2L11E,W2L12E,W2L20E,W2L21E,W2L22E;
wire W2L00F,W2L01F,W2L02F,W2L10F,W2L11F,W2L12F,W2L20F,W2L21F,W2L22F;
wire W2M000,W2M010,W2M020,W2M100,W2M110,W2M120,W2M200,W2M210,W2M220;
wire W2M001,W2M011,W2M021,W2M101,W2M111,W2M121,W2M201,W2M211,W2M221;
wire W2M002,W2M012,W2M022,W2M102,W2M112,W2M122,W2M202,W2M212,W2M222;
wire W2M003,W2M013,W2M023,W2M103,W2M113,W2M123,W2M203,W2M213,W2M223;
wire W2M004,W2M014,W2M024,W2M104,W2M114,W2M124,W2M204,W2M214,W2M224;
wire W2M005,W2M015,W2M025,W2M105,W2M115,W2M125,W2M205,W2M215,W2M225;
wire W2M006,W2M016,W2M026,W2M106,W2M116,W2M126,W2M206,W2M216,W2M226;
wire W2M007,W2M017,W2M027,W2M107,W2M117,W2M127,W2M207,W2M217,W2M227;
wire W2M008,W2M018,W2M028,W2M108,W2M118,W2M128,W2M208,W2M218,W2M228;
wire W2M009,W2M019,W2M029,W2M109,W2M119,W2M129,W2M209,W2M219,W2M229;
wire W2M00A,W2M01A,W2M02A,W2M10A,W2M11A,W2M12A,W2M20A,W2M21A,W2M22A;
wire W2M00B,W2M01B,W2M02B,W2M10B,W2M11B,W2M12B,W2M20B,W2M21B,W2M22B;
wire W2M00C,W2M01C,W2M02C,W2M10C,W2M11C,W2M12C,W2M20C,W2M21C,W2M22C;
wire W2M00D,W2M01D,W2M02D,W2M10D,W2M11D,W2M12D,W2M20D,W2M21D,W2M22D;
wire W2M00E,W2M01E,W2M02E,W2M10E,W2M11E,W2M12E,W2M20E,W2M21E,W2M22E;
wire W2M00F,W2M01F,W2M02F,W2M10F,W2M11F,W2M12F,W2M20F,W2M21F,W2M22F;
wire W2N000,W2N010,W2N020,W2N100,W2N110,W2N120,W2N200,W2N210,W2N220;
wire W2N001,W2N011,W2N021,W2N101,W2N111,W2N121,W2N201,W2N211,W2N221;
wire W2N002,W2N012,W2N022,W2N102,W2N112,W2N122,W2N202,W2N212,W2N222;
wire W2N003,W2N013,W2N023,W2N103,W2N113,W2N123,W2N203,W2N213,W2N223;
wire W2N004,W2N014,W2N024,W2N104,W2N114,W2N124,W2N204,W2N214,W2N224;
wire W2N005,W2N015,W2N025,W2N105,W2N115,W2N125,W2N205,W2N215,W2N225;
wire W2N006,W2N016,W2N026,W2N106,W2N116,W2N126,W2N206,W2N216,W2N226;
wire W2N007,W2N017,W2N027,W2N107,W2N117,W2N127,W2N207,W2N217,W2N227;
wire W2N008,W2N018,W2N028,W2N108,W2N118,W2N128,W2N208,W2N218,W2N228;
wire W2N009,W2N019,W2N029,W2N109,W2N119,W2N129,W2N209,W2N219,W2N229;
wire W2N00A,W2N01A,W2N02A,W2N10A,W2N11A,W2N12A,W2N20A,W2N21A,W2N22A;
wire W2N00B,W2N01B,W2N02B,W2N10B,W2N11B,W2N12B,W2N20B,W2N21B,W2N22B;
wire W2N00C,W2N01C,W2N02C,W2N10C,W2N11C,W2N12C,W2N20C,W2N21C,W2N22C;
wire W2N00D,W2N01D,W2N02D,W2N10D,W2N11D,W2N12D,W2N20D,W2N21D,W2N22D;
wire W2N00E,W2N01E,W2N02E,W2N10E,W2N11E,W2N12E,W2N20E,W2N21E,W2N22E;
wire W2N00F,W2N01F,W2N02F,W2N10F,W2N11F,W2N12F,W2N20F,W2N21F,W2N22F;
wire W2O000,W2O010,W2O020,W2O100,W2O110,W2O120,W2O200,W2O210,W2O220;
wire W2O001,W2O011,W2O021,W2O101,W2O111,W2O121,W2O201,W2O211,W2O221;
wire W2O002,W2O012,W2O022,W2O102,W2O112,W2O122,W2O202,W2O212,W2O222;
wire W2O003,W2O013,W2O023,W2O103,W2O113,W2O123,W2O203,W2O213,W2O223;
wire W2O004,W2O014,W2O024,W2O104,W2O114,W2O124,W2O204,W2O214,W2O224;
wire W2O005,W2O015,W2O025,W2O105,W2O115,W2O125,W2O205,W2O215,W2O225;
wire W2O006,W2O016,W2O026,W2O106,W2O116,W2O126,W2O206,W2O216,W2O226;
wire W2O007,W2O017,W2O027,W2O107,W2O117,W2O127,W2O207,W2O217,W2O227;
wire W2O008,W2O018,W2O028,W2O108,W2O118,W2O128,W2O208,W2O218,W2O228;
wire W2O009,W2O019,W2O029,W2O109,W2O119,W2O129,W2O209,W2O219,W2O229;
wire W2O00A,W2O01A,W2O02A,W2O10A,W2O11A,W2O12A,W2O20A,W2O21A,W2O22A;
wire W2O00B,W2O01B,W2O02B,W2O10B,W2O11B,W2O12B,W2O20B,W2O21B,W2O22B;
wire W2O00C,W2O01C,W2O02C,W2O10C,W2O11C,W2O12C,W2O20C,W2O21C,W2O22C;
wire W2O00D,W2O01D,W2O02D,W2O10D,W2O11D,W2O12D,W2O20D,W2O21D,W2O22D;
wire W2O00E,W2O01E,W2O02E,W2O10E,W2O11E,W2O12E,W2O20E,W2O21E,W2O22E;
wire W2O00F,W2O01F,W2O02F,W2O10F,W2O11F,W2O12F,W2O20F,W2O21F,W2O22F;
wire W2P000,W2P010,W2P020,W2P100,W2P110,W2P120,W2P200,W2P210,W2P220;
wire W2P001,W2P011,W2P021,W2P101,W2P111,W2P121,W2P201,W2P211,W2P221;
wire W2P002,W2P012,W2P022,W2P102,W2P112,W2P122,W2P202,W2P212,W2P222;
wire W2P003,W2P013,W2P023,W2P103,W2P113,W2P123,W2P203,W2P213,W2P223;
wire W2P004,W2P014,W2P024,W2P104,W2P114,W2P124,W2P204,W2P214,W2P224;
wire W2P005,W2P015,W2P025,W2P105,W2P115,W2P125,W2P205,W2P215,W2P225;
wire W2P006,W2P016,W2P026,W2P106,W2P116,W2P126,W2P206,W2P216,W2P226;
wire W2P007,W2P017,W2P027,W2P107,W2P117,W2P127,W2P207,W2P217,W2P227;
wire W2P008,W2P018,W2P028,W2P108,W2P118,W2P128,W2P208,W2P218,W2P228;
wire W2P009,W2P019,W2P029,W2P109,W2P119,W2P129,W2P209,W2P219,W2P229;
wire W2P00A,W2P01A,W2P02A,W2P10A,W2P11A,W2P12A,W2P20A,W2P21A,W2P22A;
wire W2P00B,W2P01B,W2P02B,W2P10B,W2P11B,W2P12B,W2P20B,W2P21B,W2P22B;
wire W2P00C,W2P01C,W2P02C,W2P10C,W2P11C,W2P12C,W2P20C,W2P21C,W2P22C;
wire W2P00D,W2P01D,W2P02D,W2P10D,W2P11D,W2P12D,W2P20D,W2P21D,W2P22D;
wire W2P00E,W2P01E,W2P02E,W2P10E,W2P11E,W2P12E,W2P20E,W2P21E,W2P22E;
wire W2P00F,W2P01F,W2P02F,W2P10F,W2P11F,W2P12F,W2P20F,W2P21F,W2P22F;
wire W2Q000,W2Q010,W2Q020,W2Q100,W2Q110,W2Q120,W2Q200,W2Q210,W2Q220;
wire W2Q001,W2Q011,W2Q021,W2Q101,W2Q111,W2Q121,W2Q201,W2Q211,W2Q221;
wire W2Q002,W2Q012,W2Q022,W2Q102,W2Q112,W2Q122,W2Q202,W2Q212,W2Q222;
wire W2Q003,W2Q013,W2Q023,W2Q103,W2Q113,W2Q123,W2Q203,W2Q213,W2Q223;
wire W2Q004,W2Q014,W2Q024,W2Q104,W2Q114,W2Q124,W2Q204,W2Q214,W2Q224;
wire W2Q005,W2Q015,W2Q025,W2Q105,W2Q115,W2Q125,W2Q205,W2Q215,W2Q225;
wire W2Q006,W2Q016,W2Q026,W2Q106,W2Q116,W2Q126,W2Q206,W2Q216,W2Q226;
wire W2Q007,W2Q017,W2Q027,W2Q107,W2Q117,W2Q127,W2Q207,W2Q217,W2Q227;
wire W2Q008,W2Q018,W2Q028,W2Q108,W2Q118,W2Q128,W2Q208,W2Q218,W2Q228;
wire W2Q009,W2Q019,W2Q029,W2Q109,W2Q119,W2Q129,W2Q209,W2Q219,W2Q229;
wire W2Q00A,W2Q01A,W2Q02A,W2Q10A,W2Q11A,W2Q12A,W2Q20A,W2Q21A,W2Q22A;
wire W2Q00B,W2Q01B,W2Q02B,W2Q10B,W2Q11B,W2Q12B,W2Q20B,W2Q21B,W2Q22B;
wire W2Q00C,W2Q01C,W2Q02C,W2Q10C,W2Q11C,W2Q12C,W2Q20C,W2Q21C,W2Q22C;
wire W2Q00D,W2Q01D,W2Q02D,W2Q10D,W2Q11D,W2Q12D,W2Q20D,W2Q21D,W2Q22D;
wire W2Q00E,W2Q01E,W2Q02E,W2Q10E,W2Q11E,W2Q12E,W2Q20E,W2Q21E,W2Q22E;
wire W2Q00F,W2Q01F,W2Q02F,W2Q10F,W2Q11F,W2Q12F,W2Q20F,W2Q21F,W2Q22F;
wire W2R000,W2R010,W2R020,W2R100,W2R110,W2R120,W2R200,W2R210,W2R220;
wire W2R001,W2R011,W2R021,W2R101,W2R111,W2R121,W2R201,W2R211,W2R221;
wire W2R002,W2R012,W2R022,W2R102,W2R112,W2R122,W2R202,W2R212,W2R222;
wire W2R003,W2R013,W2R023,W2R103,W2R113,W2R123,W2R203,W2R213,W2R223;
wire W2R004,W2R014,W2R024,W2R104,W2R114,W2R124,W2R204,W2R214,W2R224;
wire W2R005,W2R015,W2R025,W2R105,W2R115,W2R125,W2R205,W2R215,W2R225;
wire W2R006,W2R016,W2R026,W2R106,W2R116,W2R126,W2R206,W2R216,W2R226;
wire W2R007,W2R017,W2R027,W2R107,W2R117,W2R127,W2R207,W2R217,W2R227;
wire W2R008,W2R018,W2R028,W2R108,W2R118,W2R128,W2R208,W2R218,W2R228;
wire W2R009,W2R019,W2R029,W2R109,W2R119,W2R129,W2R209,W2R219,W2R229;
wire W2R00A,W2R01A,W2R02A,W2R10A,W2R11A,W2R12A,W2R20A,W2R21A,W2R22A;
wire W2R00B,W2R01B,W2R02B,W2R10B,W2R11B,W2R12B,W2R20B,W2R21B,W2R22B;
wire W2R00C,W2R01C,W2R02C,W2R10C,W2R11C,W2R12C,W2R20C,W2R21C,W2R22C;
wire W2R00D,W2R01D,W2R02D,W2R10D,W2R11D,W2R12D,W2R20D,W2R21D,W2R22D;
wire W2R00E,W2R01E,W2R02E,W2R10E,W2R11E,W2R12E,W2R20E,W2R21E,W2R22E;
wire W2R00F,W2R01F,W2R02F,W2R10F,W2R11F,W2R12F,W2R20F,W2R21F,W2R22F;
wire W2S000,W2S010,W2S020,W2S100,W2S110,W2S120,W2S200,W2S210,W2S220;
wire W2S001,W2S011,W2S021,W2S101,W2S111,W2S121,W2S201,W2S211,W2S221;
wire W2S002,W2S012,W2S022,W2S102,W2S112,W2S122,W2S202,W2S212,W2S222;
wire W2S003,W2S013,W2S023,W2S103,W2S113,W2S123,W2S203,W2S213,W2S223;
wire W2S004,W2S014,W2S024,W2S104,W2S114,W2S124,W2S204,W2S214,W2S224;
wire W2S005,W2S015,W2S025,W2S105,W2S115,W2S125,W2S205,W2S215,W2S225;
wire W2S006,W2S016,W2S026,W2S106,W2S116,W2S126,W2S206,W2S216,W2S226;
wire W2S007,W2S017,W2S027,W2S107,W2S117,W2S127,W2S207,W2S217,W2S227;
wire W2S008,W2S018,W2S028,W2S108,W2S118,W2S128,W2S208,W2S218,W2S228;
wire W2S009,W2S019,W2S029,W2S109,W2S119,W2S129,W2S209,W2S219,W2S229;
wire W2S00A,W2S01A,W2S02A,W2S10A,W2S11A,W2S12A,W2S20A,W2S21A,W2S22A;
wire W2S00B,W2S01B,W2S02B,W2S10B,W2S11B,W2S12B,W2S20B,W2S21B,W2S22B;
wire W2S00C,W2S01C,W2S02C,W2S10C,W2S11C,W2S12C,W2S20C,W2S21C,W2S22C;
wire W2S00D,W2S01D,W2S02D,W2S10D,W2S11D,W2S12D,W2S20D,W2S21D,W2S22D;
wire W2S00E,W2S01E,W2S02E,W2S10E,W2S11E,W2S12E,W2S20E,W2S21E,W2S22E;
wire W2S00F,W2S01F,W2S02F,W2S10F,W2S11F,W2S12F,W2S20F,W2S21F,W2S22F;
wire W2T000,W2T010,W2T020,W2T100,W2T110,W2T120,W2T200,W2T210,W2T220;
wire W2T001,W2T011,W2T021,W2T101,W2T111,W2T121,W2T201,W2T211,W2T221;
wire W2T002,W2T012,W2T022,W2T102,W2T112,W2T122,W2T202,W2T212,W2T222;
wire W2T003,W2T013,W2T023,W2T103,W2T113,W2T123,W2T203,W2T213,W2T223;
wire W2T004,W2T014,W2T024,W2T104,W2T114,W2T124,W2T204,W2T214,W2T224;
wire W2T005,W2T015,W2T025,W2T105,W2T115,W2T125,W2T205,W2T215,W2T225;
wire W2T006,W2T016,W2T026,W2T106,W2T116,W2T126,W2T206,W2T216,W2T226;
wire W2T007,W2T017,W2T027,W2T107,W2T117,W2T127,W2T207,W2T217,W2T227;
wire W2T008,W2T018,W2T028,W2T108,W2T118,W2T128,W2T208,W2T218,W2T228;
wire W2T009,W2T019,W2T029,W2T109,W2T119,W2T129,W2T209,W2T219,W2T229;
wire W2T00A,W2T01A,W2T02A,W2T10A,W2T11A,W2T12A,W2T20A,W2T21A,W2T22A;
wire W2T00B,W2T01B,W2T02B,W2T10B,W2T11B,W2T12B,W2T20B,W2T21B,W2T22B;
wire W2T00C,W2T01C,W2T02C,W2T10C,W2T11C,W2T12C,W2T20C,W2T21C,W2T22C;
wire W2T00D,W2T01D,W2T02D,W2T10D,W2T11D,W2T12D,W2T20D,W2T21D,W2T22D;
wire W2T00E,W2T01E,W2T02E,W2T10E,W2T11E,W2T12E,W2T20E,W2T21E,W2T22E;
wire W2T00F,W2T01F,W2T02F,W2T10F,W2T11F,W2T12F,W2T20F,W2T21F,W2T22F;
wire W2U000,W2U010,W2U020,W2U100,W2U110,W2U120,W2U200,W2U210,W2U220;
wire W2U001,W2U011,W2U021,W2U101,W2U111,W2U121,W2U201,W2U211,W2U221;
wire W2U002,W2U012,W2U022,W2U102,W2U112,W2U122,W2U202,W2U212,W2U222;
wire W2U003,W2U013,W2U023,W2U103,W2U113,W2U123,W2U203,W2U213,W2U223;
wire W2U004,W2U014,W2U024,W2U104,W2U114,W2U124,W2U204,W2U214,W2U224;
wire W2U005,W2U015,W2U025,W2U105,W2U115,W2U125,W2U205,W2U215,W2U225;
wire W2U006,W2U016,W2U026,W2U106,W2U116,W2U126,W2U206,W2U216,W2U226;
wire W2U007,W2U017,W2U027,W2U107,W2U117,W2U127,W2U207,W2U217,W2U227;
wire W2U008,W2U018,W2U028,W2U108,W2U118,W2U128,W2U208,W2U218,W2U228;
wire W2U009,W2U019,W2U029,W2U109,W2U119,W2U129,W2U209,W2U219,W2U229;
wire W2U00A,W2U01A,W2U02A,W2U10A,W2U11A,W2U12A,W2U20A,W2U21A,W2U22A;
wire W2U00B,W2U01B,W2U02B,W2U10B,W2U11B,W2U12B,W2U20B,W2U21B,W2U22B;
wire W2U00C,W2U01C,W2U02C,W2U10C,W2U11C,W2U12C,W2U20C,W2U21C,W2U22C;
wire W2U00D,W2U01D,W2U02D,W2U10D,W2U11D,W2U12D,W2U20D,W2U21D,W2U22D;
wire W2U00E,W2U01E,W2U02E,W2U10E,W2U11E,W2U12E,W2U20E,W2U21E,W2U22E;
wire W2U00F,W2U01F,W2U02F,W2U10F,W2U11F,W2U12F,W2U20F,W2U21F,W2U22F;
wire W2V000,W2V010,W2V020,W2V100,W2V110,W2V120,W2V200,W2V210,W2V220;
wire W2V001,W2V011,W2V021,W2V101,W2V111,W2V121,W2V201,W2V211,W2V221;
wire W2V002,W2V012,W2V022,W2V102,W2V112,W2V122,W2V202,W2V212,W2V222;
wire W2V003,W2V013,W2V023,W2V103,W2V113,W2V123,W2V203,W2V213,W2V223;
wire W2V004,W2V014,W2V024,W2V104,W2V114,W2V124,W2V204,W2V214,W2V224;
wire W2V005,W2V015,W2V025,W2V105,W2V115,W2V125,W2V205,W2V215,W2V225;
wire W2V006,W2V016,W2V026,W2V106,W2V116,W2V126,W2V206,W2V216,W2V226;
wire W2V007,W2V017,W2V027,W2V107,W2V117,W2V127,W2V207,W2V217,W2V227;
wire W2V008,W2V018,W2V028,W2V108,W2V118,W2V128,W2V208,W2V218,W2V228;
wire W2V009,W2V019,W2V029,W2V109,W2V119,W2V129,W2V209,W2V219,W2V229;
wire W2V00A,W2V01A,W2V02A,W2V10A,W2V11A,W2V12A,W2V20A,W2V21A,W2V22A;
wire W2V00B,W2V01B,W2V02B,W2V10B,W2V11B,W2V12B,W2V20B,W2V21B,W2V22B;
wire W2V00C,W2V01C,W2V02C,W2V10C,W2V11C,W2V12C,W2V20C,W2V21C,W2V22C;
wire W2V00D,W2V01D,W2V02D,W2V10D,W2V11D,W2V12D,W2V20D,W2V21D,W2V22D;
wire W2V00E,W2V01E,W2V02E,W2V10E,W2V11E,W2V12E,W2V20E,W2V21E,W2V22E;
wire W2V00F,W2V01F,W2V02F,W2V10F,W2V11F,W2V12F,W2V20F,W2V21F,W2V22F;
wire signed [4:0] c20000,c21000,c22000,c23000,c24000,c25000,c26000,c27000,c28000,c29000,c2A000,c2B000,c2C000,c2D000,c2E000,c2F000;
wire signed [4:0] c20010,c21010,c22010,c23010,c24010,c25010,c26010,c27010,c28010,c29010,c2A010,c2B010,c2C010,c2D010,c2E010,c2F010;
wire signed [4:0] c20020,c21020,c22020,c23020,c24020,c25020,c26020,c27020,c28020,c29020,c2A020,c2B020,c2C020,c2D020,c2E020,c2F020;
wire signed [4:0] c20100,c21100,c22100,c23100,c24100,c25100,c26100,c27100,c28100,c29100,c2A100,c2B100,c2C100,c2D100,c2E100,c2F100;
wire signed [4:0] c20110,c21110,c22110,c23110,c24110,c25110,c26110,c27110,c28110,c29110,c2A110,c2B110,c2C110,c2D110,c2E110,c2F110;
wire signed [4:0] c20120,c21120,c22120,c23120,c24120,c25120,c26120,c27120,c28120,c29120,c2A120,c2B120,c2C120,c2D120,c2E120,c2F120;
wire signed [4:0] c20200,c21200,c22200,c23200,c24200,c25200,c26200,c27200,c28200,c29200,c2A200,c2B200,c2C200,c2D200,c2E200,c2F200;
wire signed [4:0] c20210,c21210,c22210,c23210,c24210,c25210,c26210,c27210,c28210,c29210,c2A210,c2B210,c2C210,c2D210,c2E210,c2F210;
wire signed [4:0] c20220,c21220,c22220,c23220,c24220,c25220,c26220,c27220,c28220,c29220,c2A220,c2B220,c2C220,c2D220,c2E220,c2F220;
wire signed [4:0] c20001,c21001,c22001,c23001,c24001,c25001,c26001,c27001,c28001,c29001,c2A001,c2B001,c2C001,c2D001,c2E001,c2F001;
wire signed [4:0] c20011,c21011,c22011,c23011,c24011,c25011,c26011,c27011,c28011,c29011,c2A011,c2B011,c2C011,c2D011,c2E011,c2F011;
wire signed [4:0] c20021,c21021,c22021,c23021,c24021,c25021,c26021,c27021,c28021,c29021,c2A021,c2B021,c2C021,c2D021,c2E021,c2F021;
wire signed [4:0] c20101,c21101,c22101,c23101,c24101,c25101,c26101,c27101,c28101,c29101,c2A101,c2B101,c2C101,c2D101,c2E101,c2F101;
wire signed [4:0] c20111,c21111,c22111,c23111,c24111,c25111,c26111,c27111,c28111,c29111,c2A111,c2B111,c2C111,c2D111,c2E111,c2F111;
wire signed [4:0] c20121,c21121,c22121,c23121,c24121,c25121,c26121,c27121,c28121,c29121,c2A121,c2B121,c2C121,c2D121,c2E121,c2F121;
wire signed [4:0] c20201,c21201,c22201,c23201,c24201,c25201,c26201,c27201,c28201,c29201,c2A201,c2B201,c2C201,c2D201,c2E201,c2F201;
wire signed [4:0] c20211,c21211,c22211,c23211,c24211,c25211,c26211,c27211,c28211,c29211,c2A211,c2B211,c2C211,c2D211,c2E211,c2F211;
wire signed [4:0] c20221,c21221,c22221,c23221,c24221,c25221,c26221,c27221,c28221,c29221,c2A221,c2B221,c2C221,c2D221,c2E221,c2F221;
wire signed [4:0] c20002,c21002,c22002,c23002,c24002,c25002,c26002,c27002,c28002,c29002,c2A002,c2B002,c2C002,c2D002,c2E002,c2F002;
wire signed [4:0] c20012,c21012,c22012,c23012,c24012,c25012,c26012,c27012,c28012,c29012,c2A012,c2B012,c2C012,c2D012,c2E012,c2F012;
wire signed [4:0] c20022,c21022,c22022,c23022,c24022,c25022,c26022,c27022,c28022,c29022,c2A022,c2B022,c2C022,c2D022,c2E022,c2F022;
wire signed [4:0] c20102,c21102,c22102,c23102,c24102,c25102,c26102,c27102,c28102,c29102,c2A102,c2B102,c2C102,c2D102,c2E102,c2F102;
wire signed [4:0] c20112,c21112,c22112,c23112,c24112,c25112,c26112,c27112,c28112,c29112,c2A112,c2B112,c2C112,c2D112,c2E112,c2F112;
wire signed [4:0] c20122,c21122,c22122,c23122,c24122,c25122,c26122,c27122,c28122,c29122,c2A122,c2B122,c2C122,c2D122,c2E122,c2F122;
wire signed [4:0] c20202,c21202,c22202,c23202,c24202,c25202,c26202,c27202,c28202,c29202,c2A202,c2B202,c2C202,c2D202,c2E202,c2F202;
wire signed [4:0] c20212,c21212,c22212,c23212,c24212,c25212,c26212,c27212,c28212,c29212,c2A212,c2B212,c2C212,c2D212,c2E212,c2F212;
wire signed [4:0] c20222,c21222,c22222,c23222,c24222,c25222,c26222,c27222,c28222,c29222,c2A222,c2B222,c2C222,c2D222,c2E222,c2F222;
wire signed [4:0] c20003,c21003,c22003,c23003,c24003,c25003,c26003,c27003,c28003,c29003,c2A003,c2B003,c2C003,c2D003,c2E003,c2F003;
wire signed [4:0] c20013,c21013,c22013,c23013,c24013,c25013,c26013,c27013,c28013,c29013,c2A013,c2B013,c2C013,c2D013,c2E013,c2F013;
wire signed [4:0] c20023,c21023,c22023,c23023,c24023,c25023,c26023,c27023,c28023,c29023,c2A023,c2B023,c2C023,c2D023,c2E023,c2F023;
wire signed [4:0] c20103,c21103,c22103,c23103,c24103,c25103,c26103,c27103,c28103,c29103,c2A103,c2B103,c2C103,c2D103,c2E103,c2F103;
wire signed [4:0] c20113,c21113,c22113,c23113,c24113,c25113,c26113,c27113,c28113,c29113,c2A113,c2B113,c2C113,c2D113,c2E113,c2F113;
wire signed [4:0] c20123,c21123,c22123,c23123,c24123,c25123,c26123,c27123,c28123,c29123,c2A123,c2B123,c2C123,c2D123,c2E123,c2F123;
wire signed [4:0] c20203,c21203,c22203,c23203,c24203,c25203,c26203,c27203,c28203,c29203,c2A203,c2B203,c2C203,c2D203,c2E203,c2F203;
wire signed [4:0] c20213,c21213,c22213,c23213,c24213,c25213,c26213,c27213,c28213,c29213,c2A213,c2B213,c2C213,c2D213,c2E213,c2F213;
wire signed [4:0] c20223,c21223,c22223,c23223,c24223,c25223,c26223,c27223,c28223,c29223,c2A223,c2B223,c2C223,c2D223,c2E223,c2F223;
wire signed [4:0] c20004,c21004,c22004,c23004,c24004,c25004,c26004,c27004,c28004,c29004,c2A004,c2B004,c2C004,c2D004,c2E004,c2F004;
wire signed [4:0] c20014,c21014,c22014,c23014,c24014,c25014,c26014,c27014,c28014,c29014,c2A014,c2B014,c2C014,c2D014,c2E014,c2F014;
wire signed [4:0] c20024,c21024,c22024,c23024,c24024,c25024,c26024,c27024,c28024,c29024,c2A024,c2B024,c2C024,c2D024,c2E024,c2F024;
wire signed [4:0] c20104,c21104,c22104,c23104,c24104,c25104,c26104,c27104,c28104,c29104,c2A104,c2B104,c2C104,c2D104,c2E104,c2F104;
wire signed [4:0] c20114,c21114,c22114,c23114,c24114,c25114,c26114,c27114,c28114,c29114,c2A114,c2B114,c2C114,c2D114,c2E114,c2F114;
wire signed [4:0] c20124,c21124,c22124,c23124,c24124,c25124,c26124,c27124,c28124,c29124,c2A124,c2B124,c2C124,c2D124,c2E124,c2F124;
wire signed [4:0] c20204,c21204,c22204,c23204,c24204,c25204,c26204,c27204,c28204,c29204,c2A204,c2B204,c2C204,c2D204,c2E204,c2F204;
wire signed [4:0] c20214,c21214,c22214,c23214,c24214,c25214,c26214,c27214,c28214,c29214,c2A214,c2B214,c2C214,c2D214,c2E214,c2F214;
wire signed [4:0] c20224,c21224,c22224,c23224,c24224,c25224,c26224,c27224,c28224,c29224,c2A224,c2B224,c2C224,c2D224,c2E224,c2F224;
wire signed [4:0] c20005,c21005,c22005,c23005,c24005,c25005,c26005,c27005,c28005,c29005,c2A005,c2B005,c2C005,c2D005,c2E005,c2F005;
wire signed [4:0] c20015,c21015,c22015,c23015,c24015,c25015,c26015,c27015,c28015,c29015,c2A015,c2B015,c2C015,c2D015,c2E015,c2F015;
wire signed [4:0] c20025,c21025,c22025,c23025,c24025,c25025,c26025,c27025,c28025,c29025,c2A025,c2B025,c2C025,c2D025,c2E025,c2F025;
wire signed [4:0] c20105,c21105,c22105,c23105,c24105,c25105,c26105,c27105,c28105,c29105,c2A105,c2B105,c2C105,c2D105,c2E105,c2F105;
wire signed [4:0] c20115,c21115,c22115,c23115,c24115,c25115,c26115,c27115,c28115,c29115,c2A115,c2B115,c2C115,c2D115,c2E115,c2F115;
wire signed [4:0] c20125,c21125,c22125,c23125,c24125,c25125,c26125,c27125,c28125,c29125,c2A125,c2B125,c2C125,c2D125,c2E125,c2F125;
wire signed [4:0] c20205,c21205,c22205,c23205,c24205,c25205,c26205,c27205,c28205,c29205,c2A205,c2B205,c2C205,c2D205,c2E205,c2F205;
wire signed [4:0] c20215,c21215,c22215,c23215,c24215,c25215,c26215,c27215,c28215,c29215,c2A215,c2B215,c2C215,c2D215,c2E215,c2F215;
wire signed [4:0] c20225,c21225,c22225,c23225,c24225,c25225,c26225,c27225,c28225,c29225,c2A225,c2B225,c2C225,c2D225,c2E225,c2F225;
wire signed [4:0] c20006,c21006,c22006,c23006,c24006,c25006,c26006,c27006,c28006,c29006,c2A006,c2B006,c2C006,c2D006,c2E006,c2F006;
wire signed [4:0] c20016,c21016,c22016,c23016,c24016,c25016,c26016,c27016,c28016,c29016,c2A016,c2B016,c2C016,c2D016,c2E016,c2F016;
wire signed [4:0] c20026,c21026,c22026,c23026,c24026,c25026,c26026,c27026,c28026,c29026,c2A026,c2B026,c2C026,c2D026,c2E026,c2F026;
wire signed [4:0] c20106,c21106,c22106,c23106,c24106,c25106,c26106,c27106,c28106,c29106,c2A106,c2B106,c2C106,c2D106,c2E106,c2F106;
wire signed [4:0] c20116,c21116,c22116,c23116,c24116,c25116,c26116,c27116,c28116,c29116,c2A116,c2B116,c2C116,c2D116,c2E116,c2F116;
wire signed [4:0] c20126,c21126,c22126,c23126,c24126,c25126,c26126,c27126,c28126,c29126,c2A126,c2B126,c2C126,c2D126,c2E126,c2F126;
wire signed [4:0] c20206,c21206,c22206,c23206,c24206,c25206,c26206,c27206,c28206,c29206,c2A206,c2B206,c2C206,c2D206,c2E206,c2F206;
wire signed [4:0] c20216,c21216,c22216,c23216,c24216,c25216,c26216,c27216,c28216,c29216,c2A216,c2B216,c2C216,c2D216,c2E216,c2F216;
wire signed [4:0] c20226,c21226,c22226,c23226,c24226,c25226,c26226,c27226,c28226,c29226,c2A226,c2B226,c2C226,c2D226,c2E226,c2F226;
wire signed [4:0] c20007,c21007,c22007,c23007,c24007,c25007,c26007,c27007,c28007,c29007,c2A007,c2B007,c2C007,c2D007,c2E007,c2F007;
wire signed [4:0] c20017,c21017,c22017,c23017,c24017,c25017,c26017,c27017,c28017,c29017,c2A017,c2B017,c2C017,c2D017,c2E017,c2F017;
wire signed [4:0] c20027,c21027,c22027,c23027,c24027,c25027,c26027,c27027,c28027,c29027,c2A027,c2B027,c2C027,c2D027,c2E027,c2F027;
wire signed [4:0] c20107,c21107,c22107,c23107,c24107,c25107,c26107,c27107,c28107,c29107,c2A107,c2B107,c2C107,c2D107,c2E107,c2F107;
wire signed [4:0] c20117,c21117,c22117,c23117,c24117,c25117,c26117,c27117,c28117,c29117,c2A117,c2B117,c2C117,c2D117,c2E117,c2F117;
wire signed [4:0] c20127,c21127,c22127,c23127,c24127,c25127,c26127,c27127,c28127,c29127,c2A127,c2B127,c2C127,c2D127,c2E127,c2F127;
wire signed [4:0] c20207,c21207,c22207,c23207,c24207,c25207,c26207,c27207,c28207,c29207,c2A207,c2B207,c2C207,c2D207,c2E207,c2F207;
wire signed [4:0] c20217,c21217,c22217,c23217,c24217,c25217,c26217,c27217,c28217,c29217,c2A217,c2B217,c2C217,c2D217,c2E217,c2F217;
wire signed [4:0] c20227,c21227,c22227,c23227,c24227,c25227,c26227,c27227,c28227,c29227,c2A227,c2B227,c2C227,c2D227,c2E227,c2F227;
wire signed [4:0] c20008,c21008,c22008,c23008,c24008,c25008,c26008,c27008,c28008,c29008,c2A008,c2B008,c2C008,c2D008,c2E008,c2F008;
wire signed [4:0] c20018,c21018,c22018,c23018,c24018,c25018,c26018,c27018,c28018,c29018,c2A018,c2B018,c2C018,c2D018,c2E018,c2F018;
wire signed [4:0] c20028,c21028,c22028,c23028,c24028,c25028,c26028,c27028,c28028,c29028,c2A028,c2B028,c2C028,c2D028,c2E028,c2F028;
wire signed [4:0] c20108,c21108,c22108,c23108,c24108,c25108,c26108,c27108,c28108,c29108,c2A108,c2B108,c2C108,c2D108,c2E108,c2F108;
wire signed [4:0] c20118,c21118,c22118,c23118,c24118,c25118,c26118,c27118,c28118,c29118,c2A118,c2B118,c2C118,c2D118,c2E118,c2F118;
wire signed [4:0] c20128,c21128,c22128,c23128,c24128,c25128,c26128,c27128,c28128,c29128,c2A128,c2B128,c2C128,c2D128,c2E128,c2F128;
wire signed [4:0] c20208,c21208,c22208,c23208,c24208,c25208,c26208,c27208,c28208,c29208,c2A208,c2B208,c2C208,c2D208,c2E208,c2F208;
wire signed [4:0] c20218,c21218,c22218,c23218,c24218,c25218,c26218,c27218,c28218,c29218,c2A218,c2B218,c2C218,c2D218,c2E218,c2F218;
wire signed [4:0] c20228,c21228,c22228,c23228,c24228,c25228,c26228,c27228,c28228,c29228,c2A228,c2B228,c2C228,c2D228,c2E228,c2F228;
wire signed [4:0] c20009,c21009,c22009,c23009,c24009,c25009,c26009,c27009,c28009,c29009,c2A009,c2B009,c2C009,c2D009,c2E009,c2F009;
wire signed [4:0] c20019,c21019,c22019,c23019,c24019,c25019,c26019,c27019,c28019,c29019,c2A019,c2B019,c2C019,c2D019,c2E019,c2F019;
wire signed [4:0] c20029,c21029,c22029,c23029,c24029,c25029,c26029,c27029,c28029,c29029,c2A029,c2B029,c2C029,c2D029,c2E029,c2F029;
wire signed [4:0] c20109,c21109,c22109,c23109,c24109,c25109,c26109,c27109,c28109,c29109,c2A109,c2B109,c2C109,c2D109,c2E109,c2F109;
wire signed [4:0] c20119,c21119,c22119,c23119,c24119,c25119,c26119,c27119,c28119,c29119,c2A119,c2B119,c2C119,c2D119,c2E119,c2F119;
wire signed [4:0] c20129,c21129,c22129,c23129,c24129,c25129,c26129,c27129,c28129,c29129,c2A129,c2B129,c2C129,c2D129,c2E129,c2F129;
wire signed [4:0] c20209,c21209,c22209,c23209,c24209,c25209,c26209,c27209,c28209,c29209,c2A209,c2B209,c2C209,c2D209,c2E209,c2F209;
wire signed [4:0] c20219,c21219,c22219,c23219,c24219,c25219,c26219,c27219,c28219,c29219,c2A219,c2B219,c2C219,c2D219,c2E219,c2F219;
wire signed [4:0] c20229,c21229,c22229,c23229,c24229,c25229,c26229,c27229,c28229,c29229,c2A229,c2B229,c2C229,c2D229,c2E229,c2F229;
wire signed [4:0] c2000A,c2100A,c2200A,c2300A,c2400A,c2500A,c2600A,c2700A,c2800A,c2900A,c2A00A,c2B00A,c2C00A,c2D00A,c2E00A,c2F00A;
wire signed [4:0] c2001A,c2101A,c2201A,c2301A,c2401A,c2501A,c2601A,c2701A,c2801A,c2901A,c2A01A,c2B01A,c2C01A,c2D01A,c2E01A,c2F01A;
wire signed [4:0] c2002A,c2102A,c2202A,c2302A,c2402A,c2502A,c2602A,c2702A,c2802A,c2902A,c2A02A,c2B02A,c2C02A,c2D02A,c2E02A,c2F02A;
wire signed [4:0] c2010A,c2110A,c2210A,c2310A,c2410A,c2510A,c2610A,c2710A,c2810A,c2910A,c2A10A,c2B10A,c2C10A,c2D10A,c2E10A,c2F10A;
wire signed [4:0] c2011A,c2111A,c2211A,c2311A,c2411A,c2511A,c2611A,c2711A,c2811A,c2911A,c2A11A,c2B11A,c2C11A,c2D11A,c2E11A,c2F11A;
wire signed [4:0] c2012A,c2112A,c2212A,c2312A,c2412A,c2512A,c2612A,c2712A,c2812A,c2912A,c2A12A,c2B12A,c2C12A,c2D12A,c2E12A,c2F12A;
wire signed [4:0] c2020A,c2120A,c2220A,c2320A,c2420A,c2520A,c2620A,c2720A,c2820A,c2920A,c2A20A,c2B20A,c2C20A,c2D20A,c2E20A,c2F20A;
wire signed [4:0] c2021A,c2121A,c2221A,c2321A,c2421A,c2521A,c2621A,c2721A,c2821A,c2921A,c2A21A,c2B21A,c2C21A,c2D21A,c2E21A,c2F21A;
wire signed [4:0] c2022A,c2122A,c2222A,c2322A,c2422A,c2522A,c2622A,c2722A,c2822A,c2922A,c2A22A,c2B22A,c2C22A,c2D22A,c2E22A,c2F22A;
wire signed [4:0] c2000B,c2100B,c2200B,c2300B,c2400B,c2500B,c2600B,c2700B,c2800B,c2900B,c2A00B,c2B00B,c2C00B,c2D00B,c2E00B,c2F00B;
wire signed [4:0] c2001B,c2101B,c2201B,c2301B,c2401B,c2501B,c2601B,c2701B,c2801B,c2901B,c2A01B,c2B01B,c2C01B,c2D01B,c2E01B,c2F01B;
wire signed [4:0] c2002B,c2102B,c2202B,c2302B,c2402B,c2502B,c2602B,c2702B,c2802B,c2902B,c2A02B,c2B02B,c2C02B,c2D02B,c2E02B,c2F02B;
wire signed [4:0] c2010B,c2110B,c2210B,c2310B,c2410B,c2510B,c2610B,c2710B,c2810B,c2910B,c2A10B,c2B10B,c2C10B,c2D10B,c2E10B,c2F10B;
wire signed [4:0] c2011B,c2111B,c2211B,c2311B,c2411B,c2511B,c2611B,c2711B,c2811B,c2911B,c2A11B,c2B11B,c2C11B,c2D11B,c2E11B,c2F11B;
wire signed [4:0] c2012B,c2112B,c2212B,c2312B,c2412B,c2512B,c2612B,c2712B,c2812B,c2912B,c2A12B,c2B12B,c2C12B,c2D12B,c2E12B,c2F12B;
wire signed [4:0] c2020B,c2120B,c2220B,c2320B,c2420B,c2520B,c2620B,c2720B,c2820B,c2920B,c2A20B,c2B20B,c2C20B,c2D20B,c2E20B,c2F20B;
wire signed [4:0] c2021B,c2121B,c2221B,c2321B,c2421B,c2521B,c2621B,c2721B,c2821B,c2921B,c2A21B,c2B21B,c2C21B,c2D21B,c2E21B,c2F21B;
wire signed [4:0] c2022B,c2122B,c2222B,c2322B,c2422B,c2522B,c2622B,c2722B,c2822B,c2922B,c2A22B,c2B22B,c2C22B,c2D22B,c2E22B,c2F22B;
wire signed [4:0] c2000C,c2100C,c2200C,c2300C,c2400C,c2500C,c2600C,c2700C,c2800C,c2900C,c2A00C,c2B00C,c2C00C,c2D00C,c2E00C,c2F00C;
wire signed [4:0] c2001C,c2101C,c2201C,c2301C,c2401C,c2501C,c2601C,c2701C,c2801C,c2901C,c2A01C,c2B01C,c2C01C,c2D01C,c2E01C,c2F01C;
wire signed [4:0] c2002C,c2102C,c2202C,c2302C,c2402C,c2502C,c2602C,c2702C,c2802C,c2902C,c2A02C,c2B02C,c2C02C,c2D02C,c2E02C,c2F02C;
wire signed [4:0] c2010C,c2110C,c2210C,c2310C,c2410C,c2510C,c2610C,c2710C,c2810C,c2910C,c2A10C,c2B10C,c2C10C,c2D10C,c2E10C,c2F10C;
wire signed [4:0] c2011C,c2111C,c2211C,c2311C,c2411C,c2511C,c2611C,c2711C,c2811C,c2911C,c2A11C,c2B11C,c2C11C,c2D11C,c2E11C,c2F11C;
wire signed [4:0] c2012C,c2112C,c2212C,c2312C,c2412C,c2512C,c2612C,c2712C,c2812C,c2912C,c2A12C,c2B12C,c2C12C,c2D12C,c2E12C,c2F12C;
wire signed [4:0] c2020C,c2120C,c2220C,c2320C,c2420C,c2520C,c2620C,c2720C,c2820C,c2920C,c2A20C,c2B20C,c2C20C,c2D20C,c2E20C,c2F20C;
wire signed [4:0] c2021C,c2121C,c2221C,c2321C,c2421C,c2521C,c2621C,c2721C,c2821C,c2921C,c2A21C,c2B21C,c2C21C,c2D21C,c2E21C,c2F21C;
wire signed [4:0] c2022C,c2122C,c2222C,c2322C,c2422C,c2522C,c2622C,c2722C,c2822C,c2922C,c2A22C,c2B22C,c2C22C,c2D22C,c2E22C,c2F22C;
wire signed [4:0] c2000D,c2100D,c2200D,c2300D,c2400D,c2500D,c2600D,c2700D,c2800D,c2900D,c2A00D,c2B00D,c2C00D,c2D00D,c2E00D,c2F00D;
wire signed [4:0] c2001D,c2101D,c2201D,c2301D,c2401D,c2501D,c2601D,c2701D,c2801D,c2901D,c2A01D,c2B01D,c2C01D,c2D01D,c2E01D,c2F01D;
wire signed [4:0] c2002D,c2102D,c2202D,c2302D,c2402D,c2502D,c2602D,c2702D,c2802D,c2902D,c2A02D,c2B02D,c2C02D,c2D02D,c2E02D,c2F02D;
wire signed [4:0] c2010D,c2110D,c2210D,c2310D,c2410D,c2510D,c2610D,c2710D,c2810D,c2910D,c2A10D,c2B10D,c2C10D,c2D10D,c2E10D,c2F10D;
wire signed [4:0] c2011D,c2111D,c2211D,c2311D,c2411D,c2511D,c2611D,c2711D,c2811D,c2911D,c2A11D,c2B11D,c2C11D,c2D11D,c2E11D,c2F11D;
wire signed [4:0] c2012D,c2112D,c2212D,c2312D,c2412D,c2512D,c2612D,c2712D,c2812D,c2912D,c2A12D,c2B12D,c2C12D,c2D12D,c2E12D,c2F12D;
wire signed [4:0] c2020D,c2120D,c2220D,c2320D,c2420D,c2520D,c2620D,c2720D,c2820D,c2920D,c2A20D,c2B20D,c2C20D,c2D20D,c2E20D,c2F20D;
wire signed [4:0] c2021D,c2121D,c2221D,c2321D,c2421D,c2521D,c2621D,c2721D,c2821D,c2921D,c2A21D,c2B21D,c2C21D,c2D21D,c2E21D,c2F21D;
wire signed [4:0] c2022D,c2122D,c2222D,c2322D,c2422D,c2522D,c2622D,c2722D,c2822D,c2922D,c2A22D,c2B22D,c2C22D,c2D22D,c2E22D,c2F22D;
wire signed [4:0] c2000E,c2100E,c2200E,c2300E,c2400E,c2500E,c2600E,c2700E,c2800E,c2900E,c2A00E,c2B00E,c2C00E,c2D00E,c2E00E,c2F00E;
wire signed [4:0] c2001E,c2101E,c2201E,c2301E,c2401E,c2501E,c2601E,c2701E,c2801E,c2901E,c2A01E,c2B01E,c2C01E,c2D01E,c2E01E,c2F01E;
wire signed [4:0] c2002E,c2102E,c2202E,c2302E,c2402E,c2502E,c2602E,c2702E,c2802E,c2902E,c2A02E,c2B02E,c2C02E,c2D02E,c2E02E,c2F02E;
wire signed [4:0] c2010E,c2110E,c2210E,c2310E,c2410E,c2510E,c2610E,c2710E,c2810E,c2910E,c2A10E,c2B10E,c2C10E,c2D10E,c2E10E,c2F10E;
wire signed [4:0] c2011E,c2111E,c2211E,c2311E,c2411E,c2511E,c2611E,c2711E,c2811E,c2911E,c2A11E,c2B11E,c2C11E,c2D11E,c2E11E,c2F11E;
wire signed [4:0] c2012E,c2112E,c2212E,c2312E,c2412E,c2512E,c2612E,c2712E,c2812E,c2912E,c2A12E,c2B12E,c2C12E,c2D12E,c2E12E,c2F12E;
wire signed [4:0] c2020E,c2120E,c2220E,c2320E,c2420E,c2520E,c2620E,c2720E,c2820E,c2920E,c2A20E,c2B20E,c2C20E,c2D20E,c2E20E,c2F20E;
wire signed [4:0] c2021E,c2121E,c2221E,c2321E,c2421E,c2521E,c2621E,c2721E,c2821E,c2921E,c2A21E,c2B21E,c2C21E,c2D21E,c2E21E,c2F21E;
wire signed [4:0] c2022E,c2122E,c2222E,c2322E,c2422E,c2522E,c2622E,c2722E,c2822E,c2922E,c2A22E,c2B22E,c2C22E,c2D22E,c2E22E,c2F22E;
wire signed [4:0] c2000F,c2100F,c2200F,c2300F,c2400F,c2500F,c2600F,c2700F,c2800F,c2900F,c2A00F,c2B00F,c2C00F,c2D00F,c2E00F,c2F00F;
wire signed [4:0] c2001F,c2101F,c2201F,c2301F,c2401F,c2501F,c2601F,c2701F,c2801F,c2901F,c2A01F,c2B01F,c2C01F,c2D01F,c2E01F,c2F01F;
wire signed [4:0] c2002F,c2102F,c2202F,c2302F,c2402F,c2502F,c2602F,c2702F,c2802F,c2902F,c2A02F,c2B02F,c2C02F,c2D02F,c2E02F,c2F02F;
wire signed [4:0] c2010F,c2110F,c2210F,c2310F,c2410F,c2510F,c2610F,c2710F,c2810F,c2910F,c2A10F,c2B10F,c2C10F,c2D10F,c2E10F,c2F10F;
wire signed [4:0] c2011F,c2111F,c2211F,c2311F,c2411F,c2511F,c2611F,c2711F,c2811F,c2911F,c2A11F,c2B11F,c2C11F,c2D11F,c2E11F,c2F11F;
wire signed [4:0] c2012F,c2112F,c2212F,c2312F,c2412F,c2512F,c2612F,c2712F,c2812F,c2912F,c2A12F,c2B12F,c2C12F,c2D12F,c2E12F,c2F12F;
wire signed [4:0] c2020F,c2120F,c2220F,c2320F,c2420F,c2520F,c2620F,c2720F,c2820F,c2920F,c2A20F,c2B20F,c2C20F,c2D20F,c2E20F,c2F20F;
wire signed [4:0] c2021F,c2121F,c2221F,c2321F,c2421F,c2521F,c2621F,c2721F,c2821F,c2921F,c2A21F,c2B21F,c2C21F,c2D21F,c2E21F,c2F21F;
wire signed [4:0] c2022F,c2122F,c2222F,c2322F,c2422F,c2522F,c2622F,c2722F,c2822F,c2922F,c2A22F,c2B22F,c2C22F,c2D22F,c2E22F,c2F22F;
wire signed [4:0] c2000G,c2100G,c2200G,c2300G,c2400G,c2500G,c2600G,c2700G,c2800G,c2900G,c2A00G,c2B00G,c2C00G,c2D00G,c2E00G,c2F00G;
wire signed [4:0] c2001G,c2101G,c2201G,c2301G,c2401G,c2501G,c2601G,c2701G,c2801G,c2901G,c2A01G,c2B01G,c2C01G,c2D01G,c2E01G,c2F01G;
wire signed [4:0] c2002G,c2102G,c2202G,c2302G,c2402G,c2502G,c2602G,c2702G,c2802G,c2902G,c2A02G,c2B02G,c2C02G,c2D02G,c2E02G,c2F02G;
wire signed [4:0] c2010G,c2110G,c2210G,c2310G,c2410G,c2510G,c2610G,c2710G,c2810G,c2910G,c2A10G,c2B10G,c2C10G,c2D10G,c2E10G,c2F10G;
wire signed [4:0] c2011G,c2111G,c2211G,c2311G,c2411G,c2511G,c2611G,c2711G,c2811G,c2911G,c2A11G,c2B11G,c2C11G,c2D11G,c2E11G,c2F11G;
wire signed [4:0] c2012G,c2112G,c2212G,c2312G,c2412G,c2512G,c2612G,c2712G,c2812G,c2912G,c2A12G,c2B12G,c2C12G,c2D12G,c2E12G,c2F12G;
wire signed [4:0] c2020G,c2120G,c2220G,c2320G,c2420G,c2520G,c2620G,c2720G,c2820G,c2920G,c2A20G,c2B20G,c2C20G,c2D20G,c2E20G,c2F20G;
wire signed [4:0] c2021G,c2121G,c2221G,c2321G,c2421G,c2521G,c2621G,c2721G,c2821G,c2921G,c2A21G,c2B21G,c2C21G,c2D21G,c2E21G,c2F21G;
wire signed [4:0] c2022G,c2122G,c2222G,c2322G,c2422G,c2522G,c2622G,c2722G,c2822G,c2922G,c2A22G,c2B22G,c2C22G,c2D22G,c2E22G,c2F22G;
wire signed [4:0] c2000H,c2100H,c2200H,c2300H,c2400H,c2500H,c2600H,c2700H,c2800H,c2900H,c2A00H,c2B00H,c2C00H,c2D00H,c2E00H,c2F00H;
wire signed [4:0] c2001H,c2101H,c2201H,c2301H,c2401H,c2501H,c2601H,c2701H,c2801H,c2901H,c2A01H,c2B01H,c2C01H,c2D01H,c2E01H,c2F01H;
wire signed [4:0] c2002H,c2102H,c2202H,c2302H,c2402H,c2502H,c2602H,c2702H,c2802H,c2902H,c2A02H,c2B02H,c2C02H,c2D02H,c2E02H,c2F02H;
wire signed [4:0] c2010H,c2110H,c2210H,c2310H,c2410H,c2510H,c2610H,c2710H,c2810H,c2910H,c2A10H,c2B10H,c2C10H,c2D10H,c2E10H,c2F10H;
wire signed [4:0] c2011H,c2111H,c2211H,c2311H,c2411H,c2511H,c2611H,c2711H,c2811H,c2911H,c2A11H,c2B11H,c2C11H,c2D11H,c2E11H,c2F11H;
wire signed [4:0] c2012H,c2112H,c2212H,c2312H,c2412H,c2512H,c2612H,c2712H,c2812H,c2912H,c2A12H,c2B12H,c2C12H,c2D12H,c2E12H,c2F12H;
wire signed [4:0] c2020H,c2120H,c2220H,c2320H,c2420H,c2520H,c2620H,c2720H,c2820H,c2920H,c2A20H,c2B20H,c2C20H,c2D20H,c2E20H,c2F20H;
wire signed [4:0] c2021H,c2121H,c2221H,c2321H,c2421H,c2521H,c2621H,c2721H,c2821H,c2921H,c2A21H,c2B21H,c2C21H,c2D21H,c2E21H,c2F21H;
wire signed [4:0] c2022H,c2122H,c2222H,c2322H,c2422H,c2522H,c2622H,c2722H,c2822H,c2922H,c2A22H,c2B22H,c2C22H,c2D22H,c2E22H,c2F22H;
wire signed [4:0] c2000I,c2100I,c2200I,c2300I,c2400I,c2500I,c2600I,c2700I,c2800I,c2900I,c2A00I,c2B00I,c2C00I,c2D00I,c2E00I,c2F00I;
wire signed [4:0] c2001I,c2101I,c2201I,c2301I,c2401I,c2501I,c2601I,c2701I,c2801I,c2901I,c2A01I,c2B01I,c2C01I,c2D01I,c2E01I,c2F01I;
wire signed [4:0] c2002I,c2102I,c2202I,c2302I,c2402I,c2502I,c2602I,c2702I,c2802I,c2902I,c2A02I,c2B02I,c2C02I,c2D02I,c2E02I,c2F02I;
wire signed [4:0] c2010I,c2110I,c2210I,c2310I,c2410I,c2510I,c2610I,c2710I,c2810I,c2910I,c2A10I,c2B10I,c2C10I,c2D10I,c2E10I,c2F10I;
wire signed [4:0] c2011I,c2111I,c2211I,c2311I,c2411I,c2511I,c2611I,c2711I,c2811I,c2911I,c2A11I,c2B11I,c2C11I,c2D11I,c2E11I,c2F11I;
wire signed [4:0] c2012I,c2112I,c2212I,c2312I,c2412I,c2512I,c2612I,c2712I,c2812I,c2912I,c2A12I,c2B12I,c2C12I,c2D12I,c2E12I,c2F12I;
wire signed [4:0] c2020I,c2120I,c2220I,c2320I,c2420I,c2520I,c2620I,c2720I,c2820I,c2920I,c2A20I,c2B20I,c2C20I,c2D20I,c2E20I,c2F20I;
wire signed [4:0] c2021I,c2121I,c2221I,c2321I,c2421I,c2521I,c2621I,c2721I,c2821I,c2921I,c2A21I,c2B21I,c2C21I,c2D21I,c2E21I,c2F21I;
wire signed [4:0] c2022I,c2122I,c2222I,c2322I,c2422I,c2522I,c2622I,c2722I,c2822I,c2922I,c2A22I,c2B22I,c2C22I,c2D22I,c2E22I,c2F22I;
wire signed [4:0] c2000J,c2100J,c2200J,c2300J,c2400J,c2500J,c2600J,c2700J,c2800J,c2900J,c2A00J,c2B00J,c2C00J,c2D00J,c2E00J,c2F00J;
wire signed [4:0] c2001J,c2101J,c2201J,c2301J,c2401J,c2501J,c2601J,c2701J,c2801J,c2901J,c2A01J,c2B01J,c2C01J,c2D01J,c2E01J,c2F01J;
wire signed [4:0] c2002J,c2102J,c2202J,c2302J,c2402J,c2502J,c2602J,c2702J,c2802J,c2902J,c2A02J,c2B02J,c2C02J,c2D02J,c2E02J,c2F02J;
wire signed [4:0] c2010J,c2110J,c2210J,c2310J,c2410J,c2510J,c2610J,c2710J,c2810J,c2910J,c2A10J,c2B10J,c2C10J,c2D10J,c2E10J,c2F10J;
wire signed [4:0] c2011J,c2111J,c2211J,c2311J,c2411J,c2511J,c2611J,c2711J,c2811J,c2911J,c2A11J,c2B11J,c2C11J,c2D11J,c2E11J,c2F11J;
wire signed [4:0] c2012J,c2112J,c2212J,c2312J,c2412J,c2512J,c2612J,c2712J,c2812J,c2912J,c2A12J,c2B12J,c2C12J,c2D12J,c2E12J,c2F12J;
wire signed [4:0] c2020J,c2120J,c2220J,c2320J,c2420J,c2520J,c2620J,c2720J,c2820J,c2920J,c2A20J,c2B20J,c2C20J,c2D20J,c2E20J,c2F20J;
wire signed [4:0] c2021J,c2121J,c2221J,c2321J,c2421J,c2521J,c2621J,c2721J,c2821J,c2921J,c2A21J,c2B21J,c2C21J,c2D21J,c2E21J,c2F21J;
wire signed [4:0] c2022J,c2122J,c2222J,c2322J,c2422J,c2522J,c2622J,c2722J,c2822J,c2922J,c2A22J,c2B22J,c2C22J,c2D22J,c2E22J,c2F22J;
wire signed [4:0] c2000K,c2100K,c2200K,c2300K,c2400K,c2500K,c2600K,c2700K,c2800K,c2900K,c2A00K,c2B00K,c2C00K,c2D00K,c2E00K,c2F00K;
wire signed [4:0] c2001K,c2101K,c2201K,c2301K,c2401K,c2501K,c2601K,c2701K,c2801K,c2901K,c2A01K,c2B01K,c2C01K,c2D01K,c2E01K,c2F01K;
wire signed [4:0] c2002K,c2102K,c2202K,c2302K,c2402K,c2502K,c2602K,c2702K,c2802K,c2902K,c2A02K,c2B02K,c2C02K,c2D02K,c2E02K,c2F02K;
wire signed [4:0] c2010K,c2110K,c2210K,c2310K,c2410K,c2510K,c2610K,c2710K,c2810K,c2910K,c2A10K,c2B10K,c2C10K,c2D10K,c2E10K,c2F10K;
wire signed [4:0] c2011K,c2111K,c2211K,c2311K,c2411K,c2511K,c2611K,c2711K,c2811K,c2911K,c2A11K,c2B11K,c2C11K,c2D11K,c2E11K,c2F11K;
wire signed [4:0] c2012K,c2112K,c2212K,c2312K,c2412K,c2512K,c2612K,c2712K,c2812K,c2912K,c2A12K,c2B12K,c2C12K,c2D12K,c2E12K,c2F12K;
wire signed [4:0] c2020K,c2120K,c2220K,c2320K,c2420K,c2520K,c2620K,c2720K,c2820K,c2920K,c2A20K,c2B20K,c2C20K,c2D20K,c2E20K,c2F20K;
wire signed [4:0] c2021K,c2121K,c2221K,c2321K,c2421K,c2521K,c2621K,c2721K,c2821K,c2921K,c2A21K,c2B21K,c2C21K,c2D21K,c2E21K,c2F21K;
wire signed [4:0] c2022K,c2122K,c2222K,c2322K,c2422K,c2522K,c2622K,c2722K,c2822K,c2922K,c2A22K,c2B22K,c2C22K,c2D22K,c2E22K,c2F22K;
wire signed [4:0] c2000L,c2100L,c2200L,c2300L,c2400L,c2500L,c2600L,c2700L,c2800L,c2900L,c2A00L,c2B00L,c2C00L,c2D00L,c2E00L,c2F00L;
wire signed [4:0] c2001L,c2101L,c2201L,c2301L,c2401L,c2501L,c2601L,c2701L,c2801L,c2901L,c2A01L,c2B01L,c2C01L,c2D01L,c2E01L,c2F01L;
wire signed [4:0] c2002L,c2102L,c2202L,c2302L,c2402L,c2502L,c2602L,c2702L,c2802L,c2902L,c2A02L,c2B02L,c2C02L,c2D02L,c2E02L,c2F02L;
wire signed [4:0] c2010L,c2110L,c2210L,c2310L,c2410L,c2510L,c2610L,c2710L,c2810L,c2910L,c2A10L,c2B10L,c2C10L,c2D10L,c2E10L,c2F10L;
wire signed [4:0] c2011L,c2111L,c2211L,c2311L,c2411L,c2511L,c2611L,c2711L,c2811L,c2911L,c2A11L,c2B11L,c2C11L,c2D11L,c2E11L,c2F11L;
wire signed [4:0] c2012L,c2112L,c2212L,c2312L,c2412L,c2512L,c2612L,c2712L,c2812L,c2912L,c2A12L,c2B12L,c2C12L,c2D12L,c2E12L,c2F12L;
wire signed [4:0] c2020L,c2120L,c2220L,c2320L,c2420L,c2520L,c2620L,c2720L,c2820L,c2920L,c2A20L,c2B20L,c2C20L,c2D20L,c2E20L,c2F20L;
wire signed [4:0] c2021L,c2121L,c2221L,c2321L,c2421L,c2521L,c2621L,c2721L,c2821L,c2921L,c2A21L,c2B21L,c2C21L,c2D21L,c2E21L,c2F21L;
wire signed [4:0] c2022L,c2122L,c2222L,c2322L,c2422L,c2522L,c2622L,c2722L,c2822L,c2922L,c2A22L,c2B22L,c2C22L,c2D22L,c2E22L,c2F22L;
wire signed [4:0] c2000M,c2100M,c2200M,c2300M,c2400M,c2500M,c2600M,c2700M,c2800M,c2900M,c2A00M,c2B00M,c2C00M,c2D00M,c2E00M,c2F00M;
wire signed [4:0] c2001M,c2101M,c2201M,c2301M,c2401M,c2501M,c2601M,c2701M,c2801M,c2901M,c2A01M,c2B01M,c2C01M,c2D01M,c2E01M,c2F01M;
wire signed [4:0] c2002M,c2102M,c2202M,c2302M,c2402M,c2502M,c2602M,c2702M,c2802M,c2902M,c2A02M,c2B02M,c2C02M,c2D02M,c2E02M,c2F02M;
wire signed [4:0] c2010M,c2110M,c2210M,c2310M,c2410M,c2510M,c2610M,c2710M,c2810M,c2910M,c2A10M,c2B10M,c2C10M,c2D10M,c2E10M,c2F10M;
wire signed [4:0] c2011M,c2111M,c2211M,c2311M,c2411M,c2511M,c2611M,c2711M,c2811M,c2911M,c2A11M,c2B11M,c2C11M,c2D11M,c2E11M,c2F11M;
wire signed [4:0] c2012M,c2112M,c2212M,c2312M,c2412M,c2512M,c2612M,c2712M,c2812M,c2912M,c2A12M,c2B12M,c2C12M,c2D12M,c2E12M,c2F12M;
wire signed [4:0] c2020M,c2120M,c2220M,c2320M,c2420M,c2520M,c2620M,c2720M,c2820M,c2920M,c2A20M,c2B20M,c2C20M,c2D20M,c2E20M,c2F20M;
wire signed [4:0] c2021M,c2121M,c2221M,c2321M,c2421M,c2521M,c2621M,c2721M,c2821M,c2921M,c2A21M,c2B21M,c2C21M,c2D21M,c2E21M,c2F21M;
wire signed [4:0] c2022M,c2122M,c2222M,c2322M,c2422M,c2522M,c2622M,c2722M,c2822M,c2922M,c2A22M,c2B22M,c2C22M,c2D22M,c2E22M,c2F22M;
wire signed [4:0] c2000N,c2100N,c2200N,c2300N,c2400N,c2500N,c2600N,c2700N,c2800N,c2900N,c2A00N,c2B00N,c2C00N,c2D00N,c2E00N,c2F00N;
wire signed [4:0] c2001N,c2101N,c2201N,c2301N,c2401N,c2501N,c2601N,c2701N,c2801N,c2901N,c2A01N,c2B01N,c2C01N,c2D01N,c2E01N,c2F01N;
wire signed [4:0] c2002N,c2102N,c2202N,c2302N,c2402N,c2502N,c2602N,c2702N,c2802N,c2902N,c2A02N,c2B02N,c2C02N,c2D02N,c2E02N,c2F02N;
wire signed [4:0] c2010N,c2110N,c2210N,c2310N,c2410N,c2510N,c2610N,c2710N,c2810N,c2910N,c2A10N,c2B10N,c2C10N,c2D10N,c2E10N,c2F10N;
wire signed [4:0] c2011N,c2111N,c2211N,c2311N,c2411N,c2511N,c2611N,c2711N,c2811N,c2911N,c2A11N,c2B11N,c2C11N,c2D11N,c2E11N,c2F11N;
wire signed [4:0] c2012N,c2112N,c2212N,c2312N,c2412N,c2512N,c2612N,c2712N,c2812N,c2912N,c2A12N,c2B12N,c2C12N,c2D12N,c2E12N,c2F12N;
wire signed [4:0] c2020N,c2120N,c2220N,c2320N,c2420N,c2520N,c2620N,c2720N,c2820N,c2920N,c2A20N,c2B20N,c2C20N,c2D20N,c2E20N,c2F20N;
wire signed [4:0] c2021N,c2121N,c2221N,c2321N,c2421N,c2521N,c2621N,c2721N,c2821N,c2921N,c2A21N,c2B21N,c2C21N,c2D21N,c2E21N,c2F21N;
wire signed [4:0] c2022N,c2122N,c2222N,c2322N,c2422N,c2522N,c2622N,c2722N,c2822N,c2922N,c2A22N,c2B22N,c2C22N,c2D22N,c2E22N,c2F22N;
wire signed [4:0] c2000O,c2100O,c2200O,c2300O,c2400O,c2500O,c2600O,c2700O,c2800O,c2900O,c2A00O,c2B00O,c2C00O,c2D00O,c2E00O,c2F00O;
wire signed [4:0] c2001O,c2101O,c2201O,c2301O,c2401O,c2501O,c2601O,c2701O,c2801O,c2901O,c2A01O,c2B01O,c2C01O,c2D01O,c2E01O,c2F01O;
wire signed [4:0] c2002O,c2102O,c2202O,c2302O,c2402O,c2502O,c2602O,c2702O,c2802O,c2902O,c2A02O,c2B02O,c2C02O,c2D02O,c2E02O,c2F02O;
wire signed [4:0] c2010O,c2110O,c2210O,c2310O,c2410O,c2510O,c2610O,c2710O,c2810O,c2910O,c2A10O,c2B10O,c2C10O,c2D10O,c2E10O,c2F10O;
wire signed [4:0] c2011O,c2111O,c2211O,c2311O,c2411O,c2511O,c2611O,c2711O,c2811O,c2911O,c2A11O,c2B11O,c2C11O,c2D11O,c2E11O,c2F11O;
wire signed [4:0] c2012O,c2112O,c2212O,c2312O,c2412O,c2512O,c2612O,c2712O,c2812O,c2912O,c2A12O,c2B12O,c2C12O,c2D12O,c2E12O,c2F12O;
wire signed [4:0] c2020O,c2120O,c2220O,c2320O,c2420O,c2520O,c2620O,c2720O,c2820O,c2920O,c2A20O,c2B20O,c2C20O,c2D20O,c2E20O,c2F20O;
wire signed [4:0] c2021O,c2121O,c2221O,c2321O,c2421O,c2521O,c2621O,c2721O,c2821O,c2921O,c2A21O,c2B21O,c2C21O,c2D21O,c2E21O,c2F21O;
wire signed [4:0] c2022O,c2122O,c2222O,c2322O,c2422O,c2522O,c2622O,c2722O,c2822O,c2922O,c2A22O,c2B22O,c2C22O,c2D22O,c2E22O,c2F22O;
wire signed [4:0] c2000P,c2100P,c2200P,c2300P,c2400P,c2500P,c2600P,c2700P,c2800P,c2900P,c2A00P,c2B00P,c2C00P,c2D00P,c2E00P,c2F00P;
wire signed [4:0] c2001P,c2101P,c2201P,c2301P,c2401P,c2501P,c2601P,c2701P,c2801P,c2901P,c2A01P,c2B01P,c2C01P,c2D01P,c2E01P,c2F01P;
wire signed [4:0] c2002P,c2102P,c2202P,c2302P,c2402P,c2502P,c2602P,c2702P,c2802P,c2902P,c2A02P,c2B02P,c2C02P,c2D02P,c2E02P,c2F02P;
wire signed [4:0] c2010P,c2110P,c2210P,c2310P,c2410P,c2510P,c2610P,c2710P,c2810P,c2910P,c2A10P,c2B10P,c2C10P,c2D10P,c2E10P,c2F10P;
wire signed [4:0] c2011P,c2111P,c2211P,c2311P,c2411P,c2511P,c2611P,c2711P,c2811P,c2911P,c2A11P,c2B11P,c2C11P,c2D11P,c2E11P,c2F11P;
wire signed [4:0] c2012P,c2112P,c2212P,c2312P,c2412P,c2512P,c2612P,c2712P,c2812P,c2912P,c2A12P,c2B12P,c2C12P,c2D12P,c2E12P,c2F12P;
wire signed [4:0] c2020P,c2120P,c2220P,c2320P,c2420P,c2520P,c2620P,c2720P,c2820P,c2920P,c2A20P,c2B20P,c2C20P,c2D20P,c2E20P,c2F20P;
wire signed [4:0] c2021P,c2121P,c2221P,c2321P,c2421P,c2521P,c2621P,c2721P,c2821P,c2921P,c2A21P,c2B21P,c2C21P,c2D21P,c2E21P,c2F21P;
wire signed [4:0] c2022P,c2122P,c2222P,c2322P,c2422P,c2522P,c2622P,c2722P,c2822P,c2922P,c2A22P,c2B22P,c2C22P,c2D22P,c2E22P,c2F22P;
wire signed [4:0] c2000Q,c2100Q,c2200Q,c2300Q,c2400Q,c2500Q,c2600Q,c2700Q,c2800Q,c2900Q,c2A00Q,c2B00Q,c2C00Q,c2D00Q,c2E00Q,c2F00Q;
wire signed [4:0] c2001Q,c2101Q,c2201Q,c2301Q,c2401Q,c2501Q,c2601Q,c2701Q,c2801Q,c2901Q,c2A01Q,c2B01Q,c2C01Q,c2D01Q,c2E01Q,c2F01Q;
wire signed [4:0] c2002Q,c2102Q,c2202Q,c2302Q,c2402Q,c2502Q,c2602Q,c2702Q,c2802Q,c2902Q,c2A02Q,c2B02Q,c2C02Q,c2D02Q,c2E02Q,c2F02Q;
wire signed [4:0] c2010Q,c2110Q,c2210Q,c2310Q,c2410Q,c2510Q,c2610Q,c2710Q,c2810Q,c2910Q,c2A10Q,c2B10Q,c2C10Q,c2D10Q,c2E10Q,c2F10Q;
wire signed [4:0] c2011Q,c2111Q,c2211Q,c2311Q,c2411Q,c2511Q,c2611Q,c2711Q,c2811Q,c2911Q,c2A11Q,c2B11Q,c2C11Q,c2D11Q,c2E11Q,c2F11Q;
wire signed [4:0] c2012Q,c2112Q,c2212Q,c2312Q,c2412Q,c2512Q,c2612Q,c2712Q,c2812Q,c2912Q,c2A12Q,c2B12Q,c2C12Q,c2D12Q,c2E12Q,c2F12Q;
wire signed [4:0] c2020Q,c2120Q,c2220Q,c2320Q,c2420Q,c2520Q,c2620Q,c2720Q,c2820Q,c2920Q,c2A20Q,c2B20Q,c2C20Q,c2D20Q,c2E20Q,c2F20Q;
wire signed [4:0] c2021Q,c2121Q,c2221Q,c2321Q,c2421Q,c2521Q,c2621Q,c2721Q,c2821Q,c2921Q,c2A21Q,c2B21Q,c2C21Q,c2D21Q,c2E21Q,c2F21Q;
wire signed [4:0] c2022Q,c2122Q,c2222Q,c2322Q,c2422Q,c2522Q,c2622Q,c2722Q,c2822Q,c2922Q,c2A22Q,c2B22Q,c2C22Q,c2D22Q,c2E22Q,c2F22Q;
wire signed [4:0] c2000R,c2100R,c2200R,c2300R,c2400R,c2500R,c2600R,c2700R,c2800R,c2900R,c2A00R,c2B00R,c2C00R,c2D00R,c2E00R,c2F00R;
wire signed [4:0] c2001R,c2101R,c2201R,c2301R,c2401R,c2501R,c2601R,c2701R,c2801R,c2901R,c2A01R,c2B01R,c2C01R,c2D01R,c2E01R,c2F01R;
wire signed [4:0] c2002R,c2102R,c2202R,c2302R,c2402R,c2502R,c2602R,c2702R,c2802R,c2902R,c2A02R,c2B02R,c2C02R,c2D02R,c2E02R,c2F02R;
wire signed [4:0] c2010R,c2110R,c2210R,c2310R,c2410R,c2510R,c2610R,c2710R,c2810R,c2910R,c2A10R,c2B10R,c2C10R,c2D10R,c2E10R,c2F10R;
wire signed [4:0] c2011R,c2111R,c2211R,c2311R,c2411R,c2511R,c2611R,c2711R,c2811R,c2911R,c2A11R,c2B11R,c2C11R,c2D11R,c2E11R,c2F11R;
wire signed [4:0] c2012R,c2112R,c2212R,c2312R,c2412R,c2512R,c2612R,c2712R,c2812R,c2912R,c2A12R,c2B12R,c2C12R,c2D12R,c2E12R,c2F12R;
wire signed [4:0] c2020R,c2120R,c2220R,c2320R,c2420R,c2520R,c2620R,c2720R,c2820R,c2920R,c2A20R,c2B20R,c2C20R,c2D20R,c2E20R,c2F20R;
wire signed [4:0] c2021R,c2121R,c2221R,c2321R,c2421R,c2521R,c2621R,c2721R,c2821R,c2921R,c2A21R,c2B21R,c2C21R,c2D21R,c2E21R,c2F21R;
wire signed [4:0] c2022R,c2122R,c2222R,c2322R,c2422R,c2522R,c2622R,c2722R,c2822R,c2922R,c2A22R,c2B22R,c2C22R,c2D22R,c2E22R,c2F22R;
wire signed [4:0] c2000S,c2100S,c2200S,c2300S,c2400S,c2500S,c2600S,c2700S,c2800S,c2900S,c2A00S,c2B00S,c2C00S,c2D00S,c2E00S,c2F00S;
wire signed [4:0] c2001S,c2101S,c2201S,c2301S,c2401S,c2501S,c2601S,c2701S,c2801S,c2901S,c2A01S,c2B01S,c2C01S,c2D01S,c2E01S,c2F01S;
wire signed [4:0] c2002S,c2102S,c2202S,c2302S,c2402S,c2502S,c2602S,c2702S,c2802S,c2902S,c2A02S,c2B02S,c2C02S,c2D02S,c2E02S,c2F02S;
wire signed [4:0] c2010S,c2110S,c2210S,c2310S,c2410S,c2510S,c2610S,c2710S,c2810S,c2910S,c2A10S,c2B10S,c2C10S,c2D10S,c2E10S,c2F10S;
wire signed [4:0] c2011S,c2111S,c2211S,c2311S,c2411S,c2511S,c2611S,c2711S,c2811S,c2911S,c2A11S,c2B11S,c2C11S,c2D11S,c2E11S,c2F11S;
wire signed [4:0] c2012S,c2112S,c2212S,c2312S,c2412S,c2512S,c2612S,c2712S,c2812S,c2912S,c2A12S,c2B12S,c2C12S,c2D12S,c2E12S,c2F12S;
wire signed [4:0] c2020S,c2120S,c2220S,c2320S,c2420S,c2520S,c2620S,c2720S,c2820S,c2920S,c2A20S,c2B20S,c2C20S,c2D20S,c2E20S,c2F20S;
wire signed [4:0] c2021S,c2121S,c2221S,c2321S,c2421S,c2521S,c2621S,c2721S,c2821S,c2921S,c2A21S,c2B21S,c2C21S,c2D21S,c2E21S,c2F21S;
wire signed [4:0] c2022S,c2122S,c2222S,c2322S,c2422S,c2522S,c2622S,c2722S,c2822S,c2922S,c2A22S,c2B22S,c2C22S,c2D22S,c2E22S,c2F22S;
wire signed [4:0] c2000T,c2100T,c2200T,c2300T,c2400T,c2500T,c2600T,c2700T,c2800T,c2900T,c2A00T,c2B00T,c2C00T,c2D00T,c2E00T,c2F00T;
wire signed [4:0] c2001T,c2101T,c2201T,c2301T,c2401T,c2501T,c2601T,c2701T,c2801T,c2901T,c2A01T,c2B01T,c2C01T,c2D01T,c2E01T,c2F01T;
wire signed [4:0] c2002T,c2102T,c2202T,c2302T,c2402T,c2502T,c2602T,c2702T,c2802T,c2902T,c2A02T,c2B02T,c2C02T,c2D02T,c2E02T,c2F02T;
wire signed [4:0] c2010T,c2110T,c2210T,c2310T,c2410T,c2510T,c2610T,c2710T,c2810T,c2910T,c2A10T,c2B10T,c2C10T,c2D10T,c2E10T,c2F10T;
wire signed [4:0] c2011T,c2111T,c2211T,c2311T,c2411T,c2511T,c2611T,c2711T,c2811T,c2911T,c2A11T,c2B11T,c2C11T,c2D11T,c2E11T,c2F11T;
wire signed [4:0] c2012T,c2112T,c2212T,c2312T,c2412T,c2512T,c2612T,c2712T,c2812T,c2912T,c2A12T,c2B12T,c2C12T,c2D12T,c2E12T,c2F12T;
wire signed [4:0] c2020T,c2120T,c2220T,c2320T,c2420T,c2520T,c2620T,c2720T,c2820T,c2920T,c2A20T,c2B20T,c2C20T,c2D20T,c2E20T,c2F20T;
wire signed [4:0] c2021T,c2121T,c2221T,c2321T,c2421T,c2521T,c2621T,c2721T,c2821T,c2921T,c2A21T,c2B21T,c2C21T,c2D21T,c2E21T,c2F21T;
wire signed [4:0] c2022T,c2122T,c2222T,c2322T,c2422T,c2522T,c2622T,c2722T,c2822T,c2922T,c2A22T,c2B22T,c2C22T,c2D22T,c2E22T,c2F22T;
wire signed [4:0] c2000U,c2100U,c2200U,c2300U,c2400U,c2500U,c2600U,c2700U,c2800U,c2900U,c2A00U,c2B00U,c2C00U,c2D00U,c2E00U,c2F00U;
wire signed [4:0] c2001U,c2101U,c2201U,c2301U,c2401U,c2501U,c2601U,c2701U,c2801U,c2901U,c2A01U,c2B01U,c2C01U,c2D01U,c2E01U,c2F01U;
wire signed [4:0] c2002U,c2102U,c2202U,c2302U,c2402U,c2502U,c2602U,c2702U,c2802U,c2902U,c2A02U,c2B02U,c2C02U,c2D02U,c2E02U,c2F02U;
wire signed [4:0] c2010U,c2110U,c2210U,c2310U,c2410U,c2510U,c2610U,c2710U,c2810U,c2910U,c2A10U,c2B10U,c2C10U,c2D10U,c2E10U,c2F10U;
wire signed [4:0] c2011U,c2111U,c2211U,c2311U,c2411U,c2511U,c2611U,c2711U,c2811U,c2911U,c2A11U,c2B11U,c2C11U,c2D11U,c2E11U,c2F11U;
wire signed [4:0] c2012U,c2112U,c2212U,c2312U,c2412U,c2512U,c2612U,c2712U,c2812U,c2912U,c2A12U,c2B12U,c2C12U,c2D12U,c2E12U,c2F12U;
wire signed [4:0] c2020U,c2120U,c2220U,c2320U,c2420U,c2520U,c2620U,c2720U,c2820U,c2920U,c2A20U,c2B20U,c2C20U,c2D20U,c2E20U,c2F20U;
wire signed [4:0] c2021U,c2121U,c2221U,c2321U,c2421U,c2521U,c2621U,c2721U,c2821U,c2921U,c2A21U,c2B21U,c2C21U,c2D21U,c2E21U,c2F21U;
wire signed [4:0] c2022U,c2122U,c2222U,c2322U,c2422U,c2522U,c2622U,c2722U,c2822U,c2922U,c2A22U,c2B22U,c2C22U,c2D22U,c2E22U,c2F22U;
wire signed [4:0] c2000V,c2100V,c2200V,c2300V,c2400V,c2500V,c2600V,c2700V,c2800V,c2900V,c2A00V,c2B00V,c2C00V,c2D00V,c2E00V,c2F00V;
wire signed [4:0] c2001V,c2101V,c2201V,c2301V,c2401V,c2501V,c2601V,c2701V,c2801V,c2901V,c2A01V,c2B01V,c2C01V,c2D01V,c2E01V,c2F01V;
wire signed [4:0] c2002V,c2102V,c2202V,c2302V,c2402V,c2502V,c2602V,c2702V,c2802V,c2902V,c2A02V,c2B02V,c2C02V,c2D02V,c2E02V,c2F02V;
wire signed [4:0] c2010V,c2110V,c2210V,c2310V,c2410V,c2510V,c2610V,c2710V,c2810V,c2910V,c2A10V,c2B10V,c2C10V,c2D10V,c2E10V,c2F10V;
wire signed [4:0] c2011V,c2111V,c2211V,c2311V,c2411V,c2511V,c2611V,c2711V,c2811V,c2911V,c2A11V,c2B11V,c2C11V,c2D11V,c2E11V,c2F11V;
wire signed [4:0] c2012V,c2112V,c2212V,c2312V,c2412V,c2512V,c2612V,c2712V,c2812V,c2912V,c2A12V,c2B12V,c2C12V,c2D12V,c2E12V,c2F12V;
wire signed [4:0] c2020V,c2120V,c2220V,c2320V,c2420V,c2520V,c2620V,c2720V,c2820V,c2920V,c2A20V,c2B20V,c2C20V,c2D20V,c2E20V,c2F20V;
wire signed [4:0] c2021V,c2121V,c2221V,c2321V,c2421V,c2521V,c2621V,c2721V,c2821V,c2921V,c2A21V,c2B21V,c2C21V,c2D21V,c2E21V,c2F21V;
wire signed [4:0] c2022V,c2122V,c2222V,c2322V,c2422V,c2522V,c2622V,c2722V,c2822V,c2922V,c2A22V,c2B22V,c2C22V,c2D22V,c2E22V,c2F22V;
wire signed [9:0] C2000;
wire A2000;
wire signed [9:0] C2010;
wire A2010;
wire signed [9:0] C2020;
wire A2020;
wire signed [9:0] C2100;
wire A2100;
wire signed [9:0] C2110;
wire A2110;
wire signed [9:0] C2120;
wire A2120;
wire signed [9:0] C2200;
wire A2200;
wire signed [9:0] C2210;
wire A2210;
wire signed [9:0] C2220;
wire A2220;
wire signed [9:0] C2001;
wire A2001;
wire signed [9:0] C2011;
wire A2011;
wire signed [9:0] C2021;
wire A2021;
wire signed [9:0] C2101;
wire A2101;
wire signed [9:0] C2111;
wire A2111;
wire signed [9:0] C2121;
wire A2121;
wire signed [9:0] C2201;
wire A2201;
wire signed [9:0] C2211;
wire A2211;
wire signed [9:0] C2221;
wire A2221;
wire signed [9:0] C2002;
wire A2002;
wire signed [9:0] C2012;
wire A2012;
wire signed [9:0] C2022;
wire A2022;
wire signed [9:0] C2102;
wire A2102;
wire signed [9:0] C2112;
wire A2112;
wire signed [9:0] C2122;
wire A2122;
wire signed [9:0] C2202;
wire A2202;
wire signed [9:0] C2212;
wire A2212;
wire signed [9:0] C2222;
wire A2222;
wire signed [9:0] C2003;
wire A2003;
wire signed [9:0] C2013;
wire A2013;
wire signed [9:0] C2023;
wire A2023;
wire signed [9:0] C2103;
wire A2103;
wire signed [9:0] C2113;
wire A2113;
wire signed [9:0] C2123;
wire A2123;
wire signed [9:0] C2203;
wire A2203;
wire signed [9:0] C2213;
wire A2213;
wire signed [9:0] C2223;
wire A2223;
wire signed [9:0] C2004;
wire A2004;
wire signed [9:0] C2014;
wire A2014;
wire signed [9:0] C2024;
wire A2024;
wire signed [9:0] C2104;
wire A2104;
wire signed [9:0] C2114;
wire A2114;
wire signed [9:0] C2124;
wire A2124;
wire signed [9:0] C2204;
wire A2204;
wire signed [9:0] C2214;
wire A2214;
wire signed [9:0] C2224;
wire A2224;
wire signed [9:0] C2005;
wire A2005;
wire signed [9:0] C2015;
wire A2015;
wire signed [9:0] C2025;
wire A2025;
wire signed [9:0] C2105;
wire A2105;
wire signed [9:0] C2115;
wire A2115;
wire signed [9:0] C2125;
wire A2125;
wire signed [9:0] C2205;
wire A2205;
wire signed [9:0] C2215;
wire A2215;
wire signed [9:0] C2225;
wire A2225;
wire signed [9:0] C2006;
wire A2006;
wire signed [9:0] C2016;
wire A2016;
wire signed [9:0] C2026;
wire A2026;
wire signed [9:0] C2106;
wire A2106;
wire signed [9:0] C2116;
wire A2116;
wire signed [9:0] C2126;
wire A2126;
wire signed [9:0] C2206;
wire A2206;
wire signed [9:0] C2216;
wire A2216;
wire signed [9:0] C2226;
wire A2226;
wire signed [9:0] C2007;
wire A2007;
wire signed [9:0] C2017;
wire A2017;
wire signed [9:0] C2027;
wire A2027;
wire signed [9:0] C2107;
wire A2107;
wire signed [9:0] C2117;
wire A2117;
wire signed [9:0] C2127;
wire A2127;
wire signed [9:0] C2207;
wire A2207;
wire signed [9:0] C2217;
wire A2217;
wire signed [9:0] C2227;
wire A2227;
wire signed [9:0] C2008;
wire A2008;
wire signed [9:0] C2018;
wire A2018;
wire signed [9:0] C2028;
wire A2028;
wire signed [9:0] C2108;
wire A2108;
wire signed [9:0] C2118;
wire A2118;
wire signed [9:0] C2128;
wire A2128;
wire signed [9:0] C2208;
wire A2208;
wire signed [9:0] C2218;
wire A2218;
wire signed [9:0] C2228;
wire A2228;
wire signed [9:0] C2009;
wire A2009;
wire signed [9:0] C2019;
wire A2019;
wire signed [9:0] C2029;
wire A2029;
wire signed [9:0] C2109;
wire A2109;
wire signed [9:0] C2119;
wire A2119;
wire signed [9:0] C2129;
wire A2129;
wire signed [9:0] C2209;
wire A2209;
wire signed [9:0] C2219;
wire A2219;
wire signed [9:0] C2229;
wire A2229;
wire signed [9:0] C200A;
wire A200A;
wire signed [9:0] C201A;
wire A201A;
wire signed [9:0] C202A;
wire A202A;
wire signed [9:0] C210A;
wire A210A;
wire signed [9:0] C211A;
wire A211A;
wire signed [9:0] C212A;
wire A212A;
wire signed [9:0] C220A;
wire A220A;
wire signed [9:0] C221A;
wire A221A;
wire signed [9:0] C222A;
wire A222A;
wire signed [9:0] C200B;
wire A200B;
wire signed [9:0] C201B;
wire A201B;
wire signed [9:0] C202B;
wire A202B;
wire signed [9:0] C210B;
wire A210B;
wire signed [9:0] C211B;
wire A211B;
wire signed [9:0] C212B;
wire A212B;
wire signed [9:0] C220B;
wire A220B;
wire signed [9:0] C221B;
wire A221B;
wire signed [9:0] C222B;
wire A222B;
wire signed [9:0] C200C;
wire A200C;
wire signed [9:0] C201C;
wire A201C;
wire signed [9:0] C202C;
wire A202C;
wire signed [9:0] C210C;
wire A210C;
wire signed [9:0] C211C;
wire A211C;
wire signed [9:0] C212C;
wire A212C;
wire signed [9:0] C220C;
wire A220C;
wire signed [9:0] C221C;
wire A221C;
wire signed [9:0] C222C;
wire A222C;
wire signed [9:0] C200D;
wire A200D;
wire signed [9:0] C201D;
wire A201D;
wire signed [9:0] C202D;
wire A202D;
wire signed [9:0] C210D;
wire A210D;
wire signed [9:0] C211D;
wire A211D;
wire signed [9:0] C212D;
wire A212D;
wire signed [9:0] C220D;
wire A220D;
wire signed [9:0] C221D;
wire A221D;
wire signed [9:0] C222D;
wire A222D;
wire signed [9:0] C200E;
wire A200E;
wire signed [9:0] C201E;
wire A201E;
wire signed [9:0] C202E;
wire A202E;
wire signed [9:0] C210E;
wire A210E;
wire signed [9:0] C211E;
wire A211E;
wire signed [9:0] C212E;
wire A212E;
wire signed [9:0] C220E;
wire A220E;
wire signed [9:0] C221E;
wire A221E;
wire signed [9:0] C222E;
wire A222E;
wire signed [9:0] C200F;
wire A200F;
wire signed [9:0] C201F;
wire A201F;
wire signed [9:0] C202F;
wire A202F;
wire signed [9:0] C210F;
wire A210F;
wire signed [9:0] C211F;
wire A211F;
wire signed [9:0] C212F;
wire A212F;
wire signed [9:0] C220F;
wire A220F;
wire signed [9:0] C221F;
wire A221F;
wire signed [9:0] C222F;
wire A222F;
wire signed [9:0] C200G;
wire A200G;
wire signed [9:0] C201G;
wire A201G;
wire signed [9:0] C202G;
wire A202G;
wire signed [9:0] C210G;
wire A210G;
wire signed [9:0] C211G;
wire A211G;
wire signed [9:0] C212G;
wire A212G;
wire signed [9:0] C220G;
wire A220G;
wire signed [9:0] C221G;
wire A221G;
wire signed [9:0] C222G;
wire A222G;
wire signed [9:0] C200H;
wire A200H;
wire signed [9:0] C201H;
wire A201H;
wire signed [9:0] C202H;
wire A202H;
wire signed [9:0] C210H;
wire A210H;
wire signed [9:0] C211H;
wire A211H;
wire signed [9:0] C212H;
wire A212H;
wire signed [9:0] C220H;
wire A220H;
wire signed [9:0] C221H;
wire A221H;
wire signed [9:0] C222H;
wire A222H;
wire signed [9:0] C200I;
wire A200I;
wire signed [9:0] C201I;
wire A201I;
wire signed [9:0] C202I;
wire A202I;
wire signed [9:0] C210I;
wire A210I;
wire signed [9:0] C211I;
wire A211I;
wire signed [9:0] C212I;
wire A212I;
wire signed [9:0] C220I;
wire A220I;
wire signed [9:0] C221I;
wire A221I;
wire signed [9:0] C222I;
wire A222I;
wire signed [9:0] C200J;
wire A200J;
wire signed [9:0] C201J;
wire A201J;
wire signed [9:0] C202J;
wire A202J;
wire signed [9:0] C210J;
wire A210J;
wire signed [9:0] C211J;
wire A211J;
wire signed [9:0] C212J;
wire A212J;
wire signed [9:0] C220J;
wire A220J;
wire signed [9:0] C221J;
wire A221J;
wire signed [9:0] C222J;
wire A222J;
wire signed [9:0] C200K;
wire A200K;
wire signed [9:0] C201K;
wire A201K;
wire signed [9:0] C202K;
wire A202K;
wire signed [9:0] C210K;
wire A210K;
wire signed [9:0] C211K;
wire A211K;
wire signed [9:0] C212K;
wire A212K;
wire signed [9:0] C220K;
wire A220K;
wire signed [9:0] C221K;
wire A221K;
wire signed [9:0] C222K;
wire A222K;
wire signed [9:0] C200L;
wire A200L;
wire signed [9:0] C201L;
wire A201L;
wire signed [9:0] C202L;
wire A202L;
wire signed [9:0] C210L;
wire A210L;
wire signed [9:0] C211L;
wire A211L;
wire signed [9:0] C212L;
wire A212L;
wire signed [9:0] C220L;
wire A220L;
wire signed [9:0] C221L;
wire A221L;
wire signed [9:0] C222L;
wire A222L;
wire signed [9:0] C200M;
wire A200M;
wire signed [9:0] C201M;
wire A201M;
wire signed [9:0] C202M;
wire A202M;
wire signed [9:0] C210M;
wire A210M;
wire signed [9:0] C211M;
wire A211M;
wire signed [9:0] C212M;
wire A212M;
wire signed [9:0] C220M;
wire A220M;
wire signed [9:0] C221M;
wire A221M;
wire signed [9:0] C222M;
wire A222M;
wire signed [9:0] C200N;
wire A200N;
wire signed [9:0] C201N;
wire A201N;
wire signed [9:0] C202N;
wire A202N;
wire signed [9:0] C210N;
wire A210N;
wire signed [9:0] C211N;
wire A211N;
wire signed [9:0] C212N;
wire A212N;
wire signed [9:0] C220N;
wire A220N;
wire signed [9:0] C221N;
wire A221N;
wire signed [9:0] C222N;
wire A222N;
wire signed [9:0] C200O;
wire A200O;
wire signed [9:0] C201O;
wire A201O;
wire signed [9:0] C202O;
wire A202O;
wire signed [9:0] C210O;
wire A210O;
wire signed [9:0] C211O;
wire A211O;
wire signed [9:0] C212O;
wire A212O;
wire signed [9:0] C220O;
wire A220O;
wire signed [9:0] C221O;
wire A221O;
wire signed [9:0] C222O;
wire A222O;
wire signed [9:0] C200P;
wire A200P;
wire signed [9:0] C201P;
wire A201P;
wire signed [9:0] C202P;
wire A202P;
wire signed [9:0] C210P;
wire A210P;
wire signed [9:0] C211P;
wire A211P;
wire signed [9:0] C212P;
wire A212P;
wire signed [9:0] C220P;
wire A220P;
wire signed [9:0] C221P;
wire A221P;
wire signed [9:0] C222P;
wire A222P;
wire signed [9:0] C200Q;
wire A200Q;
wire signed [9:0] C201Q;
wire A201Q;
wire signed [9:0] C202Q;
wire A202Q;
wire signed [9:0] C210Q;
wire A210Q;
wire signed [9:0] C211Q;
wire A211Q;
wire signed [9:0] C212Q;
wire A212Q;
wire signed [9:0] C220Q;
wire A220Q;
wire signed [9:0] C221Q;
wire A221Q;
wire signed [9:0] C222Q;
wire A222Q;
wire signed [9:0] C200R;
wire A200R;
wire signed [9:0] C201R;
wire A201R;
wire signed [9:0] C202R;
wire A202R;
wire signed [9:0] C210R;
wire A210R;
wire signed [9:0] C211R;
wire A211R;
wire signed [9:0] C212R;
wire A212R;
wire signed [9:0] C220R;
wire A220R;
wire signed [9:0] C221R;
wire A221R;
wire signed [9:0] C222R;
wire A222R;
wire signed [9:0] C200S;
wire A200S;
wire signed [9:0] C201S;
wire A201S;
wire signed [9:0] C202S;
wire A202S;
wire signed [9:0] C210S;
wire A210S;
wire signed [9:0] C211S;
wire A211S;
wire signed [9:0] C212S;
wire A212S;
wire signed [9:0] C220S;
wire A220S;
wire signed [9:0] C221S;
wire A221S;
wire signed [9:0] C222S;
wire A222S;
wire signed [9:0] C200T;
wire A200T;
wire signed [9:0] C201T;
wire A201T;
wire signed [9:0] C202T;
wire A202T;
wire signed [9:0] C210T;
wire A210T;
wire signed [9:0] C211T;
wire A211T;
wire signed [9:0] C212T;
wire A212T;
wire signed [9:0] C220T;
wire A220T;
wire signed [9:0] C221T;
wire A221T;
wire signed [9:0] C222T;
wire A222T;
wire signed [9:0] C200U;
wire A200U;
wire signed [9:0] C201U;
wire A201U;
wire signed [9:0] C202U;
wire A202U;
wire signed [9:0] C210U;
wire A210U;
wire signed [9:0] C211U;
wire A211U;
wire signed [9:0] C212U;
wire A212U;
wire signed [9:0] C220U;
wire A220U;
wire signed [9:0] C221U;
wire A221U;
wire signed [9:0] C222U;
wire A222U;
wire signed [9:0] C200V;
wire A200V;
wire signed [9:0] C201V;
wire A201V;
wire signed [9:0] C202V;
wire A202V;
wire signed [9:0] C210V;
wire A210V;
wire signed [9:0] C211V;
wire A211V;
wire signed [9:0] C212V;
wire A212V;
wire signed [9:0] C220V;
wire A220V;
wire signed [9:0] C221V;
wire A221V;
wire signed [9:0] C222V;
wire A222V;
DFF_save_fm DFF_W513(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20000));
DFF_save_fm DFF_W514(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20010));
DFF_save_fm DFF_W515(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20020));
DFF_save_fm DFF_W516(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20100));
DFF_save_fm DFF_W517(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20110));
DFF_save_fm DFF_W518(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20120));
DFF_save_fm DFF_W519(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20200));
DFF_save_fm DFF_W520(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20210));
DFF_save_fm DFF_W521(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20220));
DFF_save_fm DFF_W522(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20001));
DFF_save_fm DFF_W523(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20011));
DFF_save_fm DFF_W524(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20021));
DFF_save_fm DFF_W525(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20101));
DFF_save_fm DFF_W526(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20111));
DFF_save_fm DFF_W527(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20121));
DFF_save_fm DFF_W528(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20201));
DFF_save_fm DFF_W529(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20211));
DFF_save_fm DFF_W530(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20221));
DFF_save_fm DFF_W531(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20002));
DFF_save_fm DFF_W532(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20012));
DFF_save_fm DFF_W533(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20022));
DFF_save_fm DFF_W534(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20102));
DFF_save_fm DFF_W535(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20112));
DFF_save_fm DFF_W536(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20122));
DFF_save_fm DFF_W537(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20202));
DFF_save_fm DFF_W538(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20212));
DFF_save_fm DFF_W539(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20222));
DFF_save_fm DFF_W540(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20003));
DFF_save_fm DFF_W541(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20013));
DFF_save_fm DFF_W542(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20023));
DFF_save_fm DFF_W543(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20103));
DFF_save_fm DFF_W544(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20113));
DFF_save_fm DFF_W545(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20123));
DFF_save_fm DFF_W546(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20203));
DFF_save_fm DFF_W547(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20213));
DFF_save_fm DFF_W548(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20223));
DFF_save_fm DFF_W549(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20004));
DFF_save_fm DFF_W550(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20014));
DFF_save_fm DFF_W551(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20024));
DFF_save_fm DFF_W552(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20104));
DFF_save_fm DFF_W553(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20114));
DFF_save_fm DFF_W554(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20124));
DFF_save_fm DFF_W555(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20204));
DFF_save_fm DFF_W556(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20214));
DFF_save_fm DFF_W557(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20224));
DFF_save_fm DFF_W558(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20005));
DFF_save_fm DFF_W559(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20015));
DFF_save_fm DFF_W560(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20025));
DFF_save_fm DFF_W561(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20105));
DFF_save_fm DFF_W562(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20115));
DFF_save_fm DFF_W563(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20125));
DFF_save_fm DFF_W564(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20205));
DFF_save_fm DFF_W565(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20215));
DFF_save_fm DFF_W566(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20225));
DFF_save_fm DFF_W567(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20006));
DFF_save_fm DFF_W568(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20016));
DFF_save_fm DFF_W569(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20026));
DFF_save_fm DFF_W570(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20106));
DFF_save_fm DFF_W571(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20116));
DFF_save_fm DFF_W572(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20126));
DFF_save_fm DFF_W573(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20206));
DFF_save_fm DFF_W574(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20216));
DFF_save_fm DFF_W575(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20226));
DFF_save_fm DFF_W576(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20007));
DFF_save_fm DFF_W577(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20017));
DFF_save_fm DFF_W578(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20027));
DFF_save_fm DFF_W579(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20107));
DFF_save_fm DFF_W580(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20117));
DFF_save_fm DFF_W581(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20127));
DFF_save_fm DFF_W582(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20207));
DFF_save_fm DFF_W583(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20217));
DFF_save_fm DFF_W584(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20227));
DFF_save_fm DFF_W585(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20008));
DFF_save_fm DFF_W586(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20018));
DFF_save_fm DFF_W587(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20028));
DFF_save_fm DFF_W588(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20108));
DFF_save_fm DFF_W589(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20118));
DFF_save_fm DFF_W590(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20128));
DFF_save_fm DFF_W591(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20208));
DFF_save_fm DFF_W592(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20218));
DFF_save_fm DFF_W593(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20228));
DFF_save_fm DFF_W594(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20009));
DFF_save_fm DFF_W595(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20019));
DFF_save_fm DFF_W596(.clk(clk),.rstn(rstn),.reset_value(0),.q(W20029));
DFF_save_fm DFF_W597(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20109));
DFF_save_fm DFF_W598(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20119));
DFF_save_fm DFF_W599(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20129));
DFF_save_fm DFF_W600(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20209));
DFF_save_fm DFF_W601(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20219));
DFF_save_fm DFF_W602(.clk(clk),.rstn(rstn),.reset_value(1),.q(W20229));
DFF_save_fm DFF_W603(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2000A));
DFF_save_fm DFF_W604(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2001A));
DFF_save_fm DFF_W605(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2002A));
DFF_save_fm DFF_W606(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2010A));
DFF_save_fm DFF_W607(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2011A));
DFF_save_fm DFF_W608(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2012A));
DFF_save_fm DFF_W609(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2020A));
DFF_save_fm DFF_W610(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2021A));
DFF_save_fm DFF_W611(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2022A));
DFF_save_fm DFF_W612(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2000B));
DFF_save_fm DFF_W613(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2001B));
DFF_save_fm DFF_W614(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2002B));
DFF_save_fm DFF_W615(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2010B));
DFF_save_fm DFF_W616(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2011B));
DFF_save_fm DFF_W617(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2012B));
DFF_save_fm DFF_W618(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2020B));
DFF_save_fm DFF_W619(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2021B));
DFF_save_fm DFF_W620(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2022B));
DFF_save_fm DFF_W621(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2000C));
DFF_save_fm DFF_W622(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2001C));
DFF_save_fm DFF_W623(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2002C));
DFF_save_fm DFF_W624(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2010C));
DFF_save_fm DFF_W625(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2011C));
DFF_save_fm DFF_W626(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2012C));
DFF_save_fm DFF_W627(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2020C));
DFF_save_fm DFF_W628(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2021C));
DFF_save_fm DFF_W629(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2022C));
DFF_save_fm DFF_W630(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2000D));
DFF_save_fm DFF_W631(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2001D));
DFF_save_fm DFF_W632(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2002D));
DFF_save_fm DFF_W633(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2010D));
DFF_save_fm DFF_W634(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2011D));
DFF_save_fm DFF_W635(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2012D));
DFF_save_fm DFF_W636(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2020D));
DFF_save_fm DFF_W637(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2021D));
DFF_save_fm DFF_W638(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2022D));
DFF_save_fm DFF_W639(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2000E));
DFF_save_fm DFF_W640(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2001E));
DFF_save_fm DFF_W641(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2002E));
DFF_save_fm DFF_W642(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2010E));
DFF_save_fm DFF_W643(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2011E));
DFF_save_fm DFF_W644(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2012E));
DFF_save_fm DFF_W645(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2020E));
DFF_save_fm DFF_W646(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2021E));
DFF_save_fm DFF_W647(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2022E));
DFF_save_fm DFF_W648(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2000F));
DFF_save_fm DFF_W649(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2001F));
DFF_save_fm DFF_W650(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2002F));
DFF_save_fm DFF_W651(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2010F));
DFF_save_fm DFF_W652(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2011F));
DFF_save_fm DFF_W653(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2012F));
DFF_save_fm DFF_W654(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2020F));
DFF_save_fm DFF_W655(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2021F));
DFF_save_fm DFF_W656(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2022F));
DFF_save_fm DFF_W657(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21000));
DFF_save_fm DFF_W658(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21010));
DFF_save_fm DFF_W659(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21020));
DFF_save_fm DFF_W660(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21100));
DFF_save_fm DFF_W661(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21110));
DFF_save_fm DFF_W662(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21120));
DFF_save_fm DFF_W663(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21200));
DFF_save_fm DFF_W664(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21210));
DFF_save_fm DFF_W665(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21220));
DFF_save_fm DFF_W666(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21001));
DFF_save_fm DFF_W667(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21011));
DFF_save_fm DFF_W668(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21021));
DFF_save_fm DFF_W669(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21101));
DFF_save_fm DFF_W670(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21111));
DFF_save_fm DFF_W671(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21121));
DFF_save_fm DFF_W672(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21201));
DFF_save_fm DFF_W673(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21211));
DFF_save_fm DFF_W674(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21221));
DFF_save_fm DFF_W675(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21002));
DFF_save_fm DFF_W676(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21012));
DFF_save_fm DFF_W677(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21022));
DFF_save_fm DFF_W678(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21102));
DFF_save_fm DFF_W679(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21112));
DFF_save_fm DFF_W680(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21122));
DFF_save_fm DFF_W681(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21202));
DFF_save_fm DFF_W682(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21212));
DFF_save_fm DFF_W683(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21222));
DFF_save_fm DFF_W684(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21003));
DFF_save_fm DFF_W685(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21013));
DFF_save_fm DFF_W686(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21023));
DFF_save_fm DFF_W687(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21103));
DFF_save_fm DFF_W688(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21113));
DFF_save_fm DFF_W689(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21123));
DFF_save_fm DFF_W690(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21203));
DFF_save_fm DFF_W691(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21213));
DFF_save_fm DFF_W692(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21223));
DFF_save_fm DFF_W693(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21004));
DFF_save_fm DFF_W694(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21014));
DFF_save_fm DFF_W695(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21024));
DFF_save_fm DFF_W696(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21104));
DFF_save_fm DFF_W697(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21114));
DFF_save_fm DFF_W698(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21124));
DFF_save_fm DFF_W699(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21204));
DFF_save_fm DFF_W700(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21214));
DFF_save_fm DFF_W701(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21224));
DFF_save_fm DFF_W702(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21005));
DFF_save_fm DFF_W703(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21015));
DFF_save_fm DFF_W704(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21025));
DFF_save_fm DFF_W705(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21105));
DFF_save_fm DFF_W706(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21115));
DFF_save_fm DFF_W707(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21125));
DFF_save_fm DFF_W708(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21205));
DFF_save_fm DFF_W709(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21215));
DFF_save_fm DFF_W710(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21225));
DFF_save_fm DFF_W711(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21006));
DFF_save_fm DFF_W712(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21016));
DFF_save_fm DFF_W713(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21026));
DFF_save_fm DFF_W714(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21106));
DFF_save_fm DFF_W715(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21116));
DFF_save_fm DFF_W716(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21126));
DFF_save_fm DFF_W717(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21206));
DFF_save_fm DFF_W718(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21216));
DFF_save_fm DFF_W719(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21226));
DFF_save_fm DFF_W720(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21007));
DFF_save_fm DFF_W721(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21017));
DFF_save_fm DFF_W722(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21027));
DFF_save_fm DFF_W723(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21107));
DFF_save_fm DFF_W724(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21117));
DFF_save_fm DFF_W725(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21127));
DFF_save_fm DFF_W726(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21207));
DFF_save_fm DFF_W727(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21217));
DFF_save_fm DFF_W728(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21227));
DFF_save_fm DFF_W729(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21008));
DFF_save_fm DFF_W730(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21018));
DFF_save_fm DFF_W731(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21028));
DFF_save_fm DFF_W732(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21108));
DFF_save_fm DFF_W733(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21118));
DFF_save_fm DFF_W734(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21128));
DFF_save_fm DFF_W735(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21208));
DFF_save_fm DFF_W736(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21218));
DFF_save_fm DFF_W737(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21228));
DFF_save_fm DFF_W738(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21009));
DFF_save_fm DFF_W739(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21019));
DFF_save_fm DFF_W740(.clk(clk),.rstn(rstn),.reset_value(0),.q(W21029));
DFF_save_fm DFF_W741(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21109));
DFF_save_fm DFF_W742(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21119));
DFF_save_fm DFF_W743(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21129));
DFF_save_fm DFF_W744(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21209));
DFF_save_fm DFF_W745(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21219));
DFF_save_fm DFF_W746(.clk(clk),.rstn(rstn),.reset_value(1),.q(W21229));
DFF_save_fm DFF_W747(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2100A));
DFF_save_fm DFF_W748(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2101A));
DFF_save_fm DFF_W749(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2102A));
DFF_save_fm DFF_W750(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2110A));
DFF_save_fm DFF_W751(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2111A));
DFF_save_fm DFF_W752(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2112A));
DFF_save_fm DFF_W753(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2120A));
DFF_save_fm DFF_W754(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2121A));
DFF_save_fm DFF_W755(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2122A));
DFF_save_fm DFF_W756(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2100B));
DFF_save_fm DFF_W757(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2101B));
DFF_save_fm DFF_W758(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2102B));
DFF_save_fm DFF_W759(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2110B));
DFF_save_fm DFF_W760(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2111B));
DFF_save_fm DFF_W761(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2112B));
DFF_save_fm DFF_W762(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2120B));
DFF_save_fm DFF_W763(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2121B));
DFF_save_fm DFF_W764(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2122B));
DFF_save_fm DFF_W765(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2100C));
DFF_save_fm DFF_W766(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2101C));
DFF_save_fm DFF_W767(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2102C));
DFF_save_fm DFF_W768(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2110C));
DFF_save_fm DFF_W769(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2111C));
DFF_save_fm DFF_W770(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2112C));
DFF_save_fm DFF_W771(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2120C));
DFF_save_fm DFF_W772(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2121C));
DFF_save_fm DFF_W773(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2122C));
DFF_save_fm DFF_W774(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2100D));
DFF_save_fm DFF_W775(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2101D));
DFF_save_fm DFF_W776(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2102D));
DFF_save_fm DFF_W777(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2110D));
DFF_save_fm DFF_W778(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2111D));
DFF_save_fm DFF_W779(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2112D));
DFF_save_fm DFF_W780(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2120D));
DFF_save_fm DFF_W781(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2121D));
DFF_save_fm DFF_W782(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2122D));
DFF_save_fm DFF_W783(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2100E));
DFF_save_fm DFF_W784(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2101E));
DFF_save_fm DFF_W785(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2102E));
DFF_save_fm DFF_W786(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2110E));
DFF_save_fm DFF_W787(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2111E));
DFF_save_fm DFF_W788(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2112E));
DFF_save_fm DFF_W789(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2120E));
DFF_save_fm DFF_W790(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2121E));
DFF_save_fm DFF_W791(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2122E));
DFF_save_fm DFF_W792(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2100F));
DFF_save_fm DFF_W793(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2101F));
DFF_save_fm DFF_W794(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2102F));
DFF_save_fm DFF_W795(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2110F));
DFF_save_fm DFF_W796(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2111F));
DFF_save_fm DFF_W797(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2112F));
DFF_save_fm DFF_W798(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2120F));
DFF_save_fm DFF_W799(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2121F));
DFF_save_fm DFF_W800(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2122F));
DFF_save_fm DFF_W801(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22000));
DFF_save_fm DFF_W802(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22010));
DFF_save_fm DFF_W803(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22020));
DFF_save_fm DFF_W804(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22100));
DFF_save_fm DFF_W805(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22110));
DFF_save_fm DFF_W806(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22120));
DFF_save_fm DFF_W807(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22200));
DFF_save_fm DFF_W808(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22210));
DFF_save_fm DFF_W809(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22220));
DFF_save_fm DFF_W810(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22001));
DFF_save_fm DFF_W811(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22011));
DFF_save_fm DFF_W812(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22021));
DFF_save_fm DFF_W813(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22101));
DFF_save_fm DFF_W814(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22111));
DFF_save_fm DFF_W815(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22121));
DFF_save_fm DFF_W816(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22201));
DFF_save_fm DFF_W817(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22211));
DFF_save_fm DFF_W818(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22221));
DFF_save_fm DFF_W819(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22002));
DFF_save_fm DFF_W820(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22012));
DFF_save_fm DFF_W821(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22022));
DFF_save_fm DFF_W822(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22102));
DFF_save_fm DFF_W823(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22112));
DFF_save_fm DFF_W824(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22122));
DFF_save_fm DFF_W825(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22202));
DFF_save_fm DFF_W826(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22212));
DFF_save_fm DFF_W827(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22222));
DFF_save_fm DFF_W828(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22003));
DFF_save_fm DFF_W829(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22013));
DFF_save_fm DFF_W830(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22023));
DFF_save_fm DFF_W831(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22103));
DFF_save_fm DFF_W832(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22113));
DFF_save_fm DFF_W833(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22123));
DFF_save_fm DFF_W834(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22203));
DFF_save_fm DFF_W835(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22213));
DFF_save_fm DFF_W836(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22223));
DFF_save_fm DFF_W837(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22004));
DFF_save_fm DFF_W838(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22014));
DFF_save_fm DFF_W839(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22024));
DFF_save_fm DFF_W840(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22104));
DFF_save_fm DFF_W841(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22114));
DFF_save_fm DFF_W842(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22124));
DFF_save_fm DFF_W843(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22204));
DFF_save_fm DFF_W844(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22214));
DFF_save_fm DFF_W845(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22224));
DFF_save_fm DFF_W846(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22005));
DFF_save_fm DFF_W847(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22015));
DFF_save_fm DFF_W848(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22025));
DFF_save_fm DFF_W849(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22105));
DFF_save_fm DFF_W850(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22115));
DFF_save_fm DFF_W851(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22125));
DFF_save_fm DFF_W852(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22205));
DFF_save_fm DFF_W853(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22215));
DFF_save_fm DFF_W854(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22225));
DFF_save_fm DFF_W855(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22006));
DFF_save_fm DFF_W856(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22016));
DFF_save_fm DFF_W857(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22026));
DFF_save_fm DFF_W858(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22106));
DFF_save_fm DFF_W859(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22116));
DFF_save_fm DFF_W860(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22126));
DFF_save_fm DFF_W861(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22206));
DFF_save_fm DFF_W862(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22216));
DFF_save_fm DFF_W863(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22226));
DFF_save_fm DFF_W864(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22007));
DFF_save_fm DFF_W865(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22017));
DFF_save_fm DFF_W866(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22027));
DFF_save_fm DFF_W867(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22107));
DFF_save_fm DFF_W868(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22117));
DFF_save_fm DFF_W869(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22127));
DFF_save_fm DFF_W870(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22207));
DFF_save_fm DFF_W871(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22217));
DFF_save_fm DFF_W872(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22227));
DFF_save_fm DFF_W873(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22008));
DFF_save_fm DFF_W874(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22018));
DFF_save_fm DFF_W875(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22028));
DFF_save_fm DFF_W876(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22108));
DFF_save_fm DFF_W877(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22118));
DFF_save_fm DFF_W878(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22128));
DFF_save_fm DFF_W879(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22208));
DFF_save_fm DFF_W880(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22218));
DFF_save_fm DFF_W881(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22228));
DFF_save_fm DFF_W882(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22009));
DFF_save_fm DFF_W883(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22019));
DFF_save_fm DFF_W884(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22029));
DFF_save_fm DFF_W885(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22109));
DFF_save_fm DFF_W886(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22119));
DFF_save_fm DFF_W887(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22129));
DFF_save_fm DFF_W888(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22209));
DFF_save_fm DFF_W889(.clk(clk),.rstn(rstn),.reset_value(1),.q(W22219));
DFF_save_fm DFF_W890(.clk(clk),.rstn(rstn),.reset_value(0),.q(W22229));
DFF_save_fm DFF_W891(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2200A));
DFF_save_fm DFF_W892(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2201A));
DFF_save_fm DFF_W893(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2202A));
DFF_save_fm DFF_W894(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2210A));
DFF_save_fm DFF_W895(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2211A));
DFF_save_fm DFF_W896(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2212A));
DFF_save_fm DFF_W897(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2220A));
DFF_save_fm DFF_W898(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2221A));
DFF_save_fm DFF_W899(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2222A));
DFF_save_fm DFF_W900(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2200B));
DFF_save_fm DFF_W901(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2201B));
DFF_save_fm DFF_W902(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2202B));
DFF_save_fm DFF_W903(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2210B));
DFF_save_fm DFF_W904(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2211B));
DFF_save_fm DFF_W905(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2212B));
DFF_save_fm DFF_W906(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2220B));
DFF_save_fm DFF_W907(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2221B));
DFF_save_fm DFF_W908(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2222B));
DFF_save_fm DFF_W909(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2200C));
DFF_save_fm DFF_W910(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2201C));
DFF_save_fm DFF_W911(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2202C));
DFF_save_fm DFF_W912(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2210C));
DFF_save_fm DFF_W913(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2211C));
DFF_save_fm DFF_W914(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2212C));
DFF_save_fm DFF_W915(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2220C));
DFF_save_fm DFF_W916(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2221C));
DFF_save_fm DFF_W917(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2222C));
DFF_save_fm DFF_W918(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2200D));
DFF_save_fm DFF_W919(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2201D));
DFF_save_fm DFF_W920(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2202D));
DFF_save_fm DFF_W921(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2210D));
DFF_save_fm DFF_W922(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2211D));
DFF_save_fm DFF_W923(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2212D));
DFF_save_fm DFF_W924(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2220D));
DFF_save_fm DFF_W925(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2221D));
DFF_save_fm DFF_W926(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2222D));
DFF_save_fm DFF_W927(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2200E));
DFF_save_fm DFF_W928(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2201E));
DFF_save_fm DFF_W929(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2202E));
DFF_save_fm DFF_W930(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2210E));
DFF_save_fm DFF_W931(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2211E));
DFF_save_fm DFF_W932(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2212E));
DFF_save_fm DFF_W933(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2220E));
DFF_save_fm DFF_W934(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2221E));
DFF_save_fm DFF_W935(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2222E));
DFF_save_fm DFF_W936(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2200F));
DFF_save_fm DFF_W937(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2201F));
DFF_save_fm DFF_W938(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2202F));
DFF_save_fm DFF_W939(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2210F));
DFF_save_fm DFF_W940(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2211F));
DFF_save_fm DFF_W941(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2212F));
DFF_save_fm DFF_W942(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2220F));
DFF_save_fm DFF_W943(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2221F));
DFF_save_fm DFF_W944(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2222F));
DFF_save_fm DFF_W945(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23000));
DFF_save_fm DFF_W946(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23010));
DFF_save_fm DFF_W947(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23020));
DFF_save_fm DFF_W948(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23100));
DFF_save_fm DFF_W949(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23110));
DFF_save_fm DFF_W950(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23120));
DFF_save_fm DFF_W951(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23200));
DFF_save_fm DFF_W952(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23210));
DFF_save_fm DFF_W953(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23220));
DFF_save_fm DFF_W954(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23001));
DFF_save_fm DFF_W955(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23011));
DFF_save_fm DFF_W956(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23021));
DFF_save_fm DFF_W957(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23101));
DFF_save_fm DFF_W958(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23111));
DFF_save_fm DFF_W959(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23121));
DFF_save_fm DFF_W960(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23201));
DFF_save_fm DFF_W961(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23211));
DFF_save_fm DFF_W962(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23221));
DFF_save_fm DFF_W963(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23002));
DFF_save_fm DFF_W964(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23012));
DFF_save_fm DFF_W965(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23022));
DFF_save_fm DFF_W966(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23102));
DFF_save_fm DFF_W967(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23112));
DFF_save_fm DFF_W968(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23122));
DFF_save_fm DFF_W969(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23202));
DFF_save_fm DFF_W970(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23212));
DFF_save_fm DFF_W971(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23222));
DFF_save_fm DFF_W972(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23003));
DFF_save_fm DFF_W973(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23013));
DFF_save_fm DFF_W974(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23023));
DFF_save_fm DFF_W975(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23103));
DFF_save_fm DFF_W976(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23113));
DFF_save_fm DFF_W977(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23123));
DFF_save_fm DFF_W978(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23203));
DFF_save_fm DFF_W979(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23213));
DFF_save_fm DFF_W980(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23223));
DFF_save_fm DFF_W981(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23004));
DFF_save_fm DFF_W982(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23014));
DFF_save_fm DFF_W983(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23024));
DFF_save_fm DFF_W984(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23104));
DFF_save_fm DFF_W985(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23114));
DFF_save_fm DFF_W986(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23124));
DFF_save_fm DFF_W987(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23204));
DFF_save_fm DFF_W988(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23214));
DFF_save_fm DFF_W989(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23224));
DFF_save_fm DFF_W990(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23005));
DFF_save_fm DFF_W991(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23015));
DFF_save_fm DFF_W992(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23025));
DFF_save_fm DFF_W993(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23105));
DFF_save_fm DFF_W994(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23115));
DFF_save_fm DFF_W995(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23125));
DFF_save_fm DFF_W996(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23205));
DFF_save_fm DFF_W997(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23215));
DFF_save_fm DFF_W998(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23225));
DFF_save_fm DFF_W999(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23006));
DFF_save_fm DFF_W1000(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23016));
DFF_save_fm DFF_W1001(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23026));
DFF_save_fm DFF_W1002(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23106));
DFF_save_fm DFF_W1003(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23116));
DFF_save_fm DFF_W1004(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23126));
DFF_save_fm DFF_W1005(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23206));
DFF_save_fm DFF_W1006(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23216));
DFF_save_fm DFF_W1007(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23226));
DFF_save_fm DFF_W1008(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23007));
DFF_save_fm DFF_W1009(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23017));
DFF_save_fm DFF_W1010(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23027));
DFF_save_fm DFF_W1011(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23107));
DFF_save_fm DFF_W1012(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23117));
DFF_save_fm DFF_W1013(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23127));
DFF_save_fm DFF_W1014(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23207));
DFF_save_fm DFF_W1015(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23217));
DFF_save_fm DFF_W1016(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23227));
DFF_save_fm DFF_W1017(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23008));
DFF_save_fm DFF_W1018(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23018));
DFF_save_fm DFF_W1019(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23028));
DFF_save_fm DFF_W1020(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23108));
DFF_save_fm DFF_W1021(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23118));
DFF_save_fm DFF_W1022(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23128));
DFF_save_fm DFF_W1023(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23208));
DFF_save_fm DFF_W1024(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23218));
DFF_save_fm DFF_W1025(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23228));
DFF_save_fm DFF_W1026(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23009));
DFF_save_fm DFF_W1027(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23019));
DFF_save_fm DFF_W1028(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23029));
DFF_save_fm DFF_W1029(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23109));
DFF_save_fm DFF_W1030(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23119));
DFF_save_fm DFF_W1031(.clk(clk),.rstn(rstn),.reset_value(0),.q(W23129));
DFF_save_fm DFF_W1032(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23209));
DFF_save_fm DFF_W1033(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23219));
DFF_save_fm DFF_W1034(.clk(clk),.rstn(rstn),.reset_value(1),.q(W23229));
DFF_save_fm DFF_W1035(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2300A));
DFF_save_fm DFF_W1036(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2301A));
DFF_save_fm DFF_W1037(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2302A));
DFF_save_fm DFF_W1038(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2310A));
DFF_save_fm DFF_W1039(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2311A));
DFF_save_fm DFF_W1040(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2312A));
DFF_save_fm DFF_W1041(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2320A));
DFF_save_fm DFF_W1042(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2321A));
DFF_save_fm DFF_W1043(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2322A));
DFF_save_fm DFF_W1044(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2300B));
DFF_save_fm DFF_W1045(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2301B));
DFF_save_fm DFF_W1046(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2302B));
DFF_save_fm DFF_W1047(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2310B));
DFF_save_fm DFF_W1048(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2311B));
DFF_save_fm DFF_W1049(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2312B));
DFF_save_fm DFF_W1050(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2320B));
DFF_save_fm DFF_W1051(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2321B));
DFF_save_fm DFF_W1052(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2322B));
DFF_save_fm DFF_W1053(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2300C));
DFF_save_fm DFF_W1054(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2301C));
DFF_save_fm DFF_W1055(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2302C));
DFF_save_fm DFF_W1056(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2310C));
DFF_save_fm DFF_W1057(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2311C));
DFF_save_fm DFF_W1058(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2312C));
DFF_save_fm DFF_W1059(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2320C));
DFF_save_fm DFF_W1060(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2321C));
DFF_save_fm DFF_W1061(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2322C));
DFF_save_fm DFF_W1062(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2300D));
DFF_save_fm DFF_W1063(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2301D));
DFF_save_fm DFF_W1064(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2302D));
DFF_save_fm DFF_W1065(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2310D));
DFF_save_fm DFF_W1066(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2311D));
DFF_save_fm DFF_W1067(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2312D));
DFF_save_fm DFF_W1068(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2320D));
DFF_save_fm DFF_W1069(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2321D));
DFF_save_fm DFF_W1070(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2322D));
DFF_save_fm DFF_W1071(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2300E));
DFF_save_fm DFF_W1072(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2301E));
DFF_save_fm DFF_W1073(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2302E));
DFF_save_fm DFF_W1074(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2310E));
DFF_save_fm DFF_W1075(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2311E));
DFF_save_fm DFF_W1076(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2312E));
DFF_save_fm DFF_W1077(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2320E));
DFF_save_fm DFF_W1078(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2321E));
DFF_save_fm DFF_W1079(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2322E));
DFF_save_fm DFF_W1080(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2300F));
DFF_save_fm DFF_W1081(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2301F));
DFF_save_fm DFF_W1082(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2302F));
DFF_save_fm DFF_W1083(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2310F));
DFF_save_fm DFF_W1084(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2311F));
DFF_save_fm DFF_W1085(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2312F));
DFF_save_fm DFF_W1086(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2320F));
DFF_save_fm DFF_W1087(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2321F));
DFF_save_fm DFF_W1088(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2322F));
DFF_save_fm DFF_W1089(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24000));
DFF_save_fm DFF_W1090(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24010));
DFF_save_fm DFF_W1091(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24020));
DFF_save_fm DFF_W1092(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24100));
DFF_save_fm DFF_W1093(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24110));
DFF_save_fm DFF_W1094(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24120));
DFF_save_fm DFF_W1095(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24200));
DFF_save_fm DFF_W1096(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24210));
DFF_save_fm DFF_W1097(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24220));
DFF_save_fm DFF_W1098(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24001));
DFF_save_fm DFF_W1099(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24011));
DFF_save_fm DFF_W1100(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24021));
DFF_save_fm DFF_W1101(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24101));
DFF_save_fm DFF_W1102(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24111));
DFF_save_fm DFF_W1103(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24121));
DFF_save_fm DFF_W1104(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24201));
DFF_save_fm DFF_W1105(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24211));
DFF_save_fm DFF_W1106(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24221));
DFF_save_fm DFF_W1107(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24002));
DFF_save_fm DFF_W1108(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24012));
DFF_save_fm DFF_W1109(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24022));
DFF_save_fm DFF_W1110(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24102));
DFF_save_fm DFF_W1111(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24112));
DFF_save_fm DFF_W1112(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24122));
DFF_save_fm DFF_W1113(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24202));
DFF_save_fm DFF_W1114(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24212));
DFF_save_fm DFF_W1115(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24222));
DFF_save_fm DFF_W1116(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24003));
DFF_save_fm DFF_W1117(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24013));
DFF_save_fm DFF_W1118(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24023));
DFF_save_fm DFF_W1119(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24103));
DFF_save_fm DFF_W1120(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24113));
DFF_save_fm DFF_W1121(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24123));
DFF_save_fm DFF_W1122(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24203));
DFF_save_fm DFF_W1123(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24213));
DFF_save_fm DFF_W1124(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24223));
DFF_save_fm DFF_W1125(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24004));
DFF_save_fm DFF_W1126(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24014));
DFF_save_fm DFF_W1127(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24024));
DFF_save_fm DFF_W1128(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24104));
DFF_save_fm DFF_W1129(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24114));
DFF_save_fm DFF_W1130(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24124));
DFF_save_fm DFF_W1131(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24204));
DFF_save_fm DFF_W1132(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24214));
DFF_save_fm DFF_W1133(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24224));
DFF_save_fm DFF_W1134(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24005));
DFF_save_fm DFF_W1135(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24015));
DFF_save_fm DFF_W1136(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24025));
DFF_save_fm DFF_W1137(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24105));
DFF_save_fm DFF_W1138(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24115));
DFF_save_fm DFF_W1139(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24125));
DFF_save_fm DFF_W1140(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24205));
DFF_save_fm DFF_W1141(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24215));
DFF_save_fm DFF_W1142(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24225));
DFF_save_fm DFF_W1143(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24006));
DFF_save_fm DFF_W1144(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24016));
DFF_save_fm DFF_W1145(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24026));
DFF_save_fm DFF_W1146(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24106));
DFF_save_fm DFF_W1147(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24116));
DFF_save_fm DFF_W1148(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24126));
DFF_save_fm DFF_W1149(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24206));
DFF_save_fm DFF_W1150(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24216));
DFF_save_fm DFF_W1151(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24226));
DFF_save_fm DFF_W1152(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24007));
DFF_save_fm DFF_W1153(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24017));
DFF_save_fm DFF_W1154(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24027));
DFF_save_fm DFF_W1155(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24107));
DFF_save_fm DFF_W1156(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24117));
DFF_save_fm DFF_W1157(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24127));
DFF_save_fm DFF_W1158(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24207));
DFF_save_fm DFF_W1159(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24217));
DFF_save_fm DFF_W1160(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24227));
DFF_save_fm DFF_W1161(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24008));
DFF_save_fm DFF_W1162(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24018));
DFF_save_fm DFF_W1163(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24028));
DFF_save_fm DFF_W1164(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24108));
DFF_save_fm DFF_W1165(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24118));
DFF_save_fm DFF_W1166(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24128));
DFF_save_fm DFF_W1167(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24208));
DFF_save_fm DFF_W1168(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24218));
DFF_save_fm DFF_W1169(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24228));
DFF_save_fm DFF_W1170(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24009));
DFF_save_fm DFF_W1171(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24019));
DFF_save_fm DFF_W1172(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24029));
DFF_save_fm DFF_W1173(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24109));
DFF_save_fm DFF_W1174(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24119));
DFF_save_fm DFF_W1175(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24129));
DFF_save_fm DFF_W1176(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24209));
DFF_save_fm DFF_W1177(.clk(clk),.rstn(rstn),.reset_value(1),.q(W24219));
DFF_save_fm DFF_W1178(.clk(clk),.rstn(rstn),.reset_value(0),.q(W24229));
DFF_save_fm DFF_W1179(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2400A));
DFF_save_fm DFF_W1180(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2401A));
DFF_save_fm DFF_W1181(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2402A));
DFF_save_fm DFF_W1182(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2410A));
DFF_save_fm DFF_W1183(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2411A));
DFF_save_fm DFF_W1184(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2412A));
DFF_save_fm DFF_W1185(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2420A));
DFF_save_fm DFF_W1186(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2421A));
DFF_save_fm DFF_W1187(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2422A));
DFF_save_fm DFF_W1188(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2400B));
DFF_save_fm DFF_W1189(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2401B));
DFF_save_fm DFF_W1190(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2402B));
DFF_save_fm DFF_W1191(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2410B));
DFF_save_fm DFF_W1192(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2411B));
DFF_save_fm DFF_W1193(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2412B));
DFF_save_fm DFF_W1194(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2420B));
DFF_save_fm DFF_W1195(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2421B));
DFF_save_fm DFF_W1196(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2422B));
DFF_save_fm DFF_W1197(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2400C));
DFF_save_fm DFF_W1198(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2401C));
DFF_save_fm DFF_W1199(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2402C));
DFF_save_fm DFF_W1200(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2410C));
DFF_save_fm DFF_W1201(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2411C));
DFF_save_fm DFF_W1202(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2412C));
DFF_save_fm DFF_W1203(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2420C));
DFF_save_fm DFF_W1204(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2421C));
DFF_save_fm DFF_W1205(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2422C));
DFF_save_fm DFF_W1206(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2400D));
DFF_save_fm DFF_W1207(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2401D));
DFF_save_fm DFF_W1208(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2402D));
DFF_save_fm DFF_W1209(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2410D));
DFF_save_fm DFF_W1210(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2411D));
DFF_save_fm DFF_W1211(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2412D));
DFF_save_fm DFF_W1212(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2420D));
DFF_save_fm DFF_W1213(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2421D));
DFF_save_fm DFF_W1214(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2422D));
DFF_save_fm DFF_W1215(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2400E));
DFF_save_fm DFF_W1216(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2401E));
DFF_save_fm DFF_W1217(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2402E));
DFF_save_fm DFF_W1218(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2410E));
DFF_save_fm DFF_W1219(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2411E));
DFF_save_fm DFF_W1220(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2412E));
DFF_save_fm DFF_W1221(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2420E));
DFF_save_fm DFF_W1222(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2421E));
DFF_save_fm DFF_W1223(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2422E));
DFF_save_fm DFF_W1224(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2400F));
DFF_save_fm DFF_W1225(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2401F));
DFF_save_fm DFF_W1226(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2402F));
DFF_save_fm DFF_W1227(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2410F));
DFF_save_fm DFF_W1228(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2411F));
DFF_save_fm DFF_W1229(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2412F));
DFF_save_fm DFF_W1230(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2420F));
DFF_save_fm DFF_W1231(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2421F));
DFF_save_fm DFF_W1232(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2422F));
DFF_save_fm DFF_W1233(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25000));
DFF_save_fm DFF_W1234(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25010));
DFF_save_fm DFF_W1235(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25020));
DFF_save_fm DFF_W1236(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25100));
DFF_save_fm DFF_W1237(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25110));
DFF_save_fm DFF_W1238(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25120));
DFF_save_fm DFF_W1239(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25200));
DFF_save_fm DFF_W1240(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25210));
DFF_save_fm DFF_W1241(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25220));
DFF_save_fm DFF_W1242(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25001));
DFF_save_fm DFF_W1243(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25011));
DFF_save_fm DFF_W1244(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25021));
DFF_save_fm DFF_W1245(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25101));
DFF_save_fm DFF_W1246(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25111));
DFF_save_fm DFF_W1247(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25121));
DFF_save_fm DFF_W1248(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25201));
DFF_save_fm DFF_W1249(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25211));
DFF_save_fm DFF_W1250(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25221));
DFF_save_fm DFF_W1251(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25002));
DFF_save_fm DFF_W1252(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25012));
DFF_save_fm DFF_W1253(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25022));
DFF_save_fm DFF_W1254(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25102));
DFF_save_fm DFF_W1255(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25112));
DFF_save_fm DFF_W1256(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25122));
DFF_save_fm DFF_W1257(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25202));
DFF_save_fm DFF_W1258(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25212));
DFF_save_fm DFF_W1259(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25222));
DFF_save_fm DFF_W1260(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25003));
DFF_save_fm DFF_W1261(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25013));
DFF_save_fm DFF_W1262(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25023));
DFF_save_fm DFF_W1263(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25103));
DFF_save_fm DFF_W1264(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25113));
DFF_save_fm DFF_W1265(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25123));
DFF_save_fm DFF_W1266(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25203));
DFF_save_fm DFF_W1267(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25213));
DFF_save_fm DFF_W1268(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25223));
DFF_save_fm DFF_W1269(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25004));
DFF_save_fm DFF_W1270(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25014));
DFF_save_fm DFF_W1271(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25024));
DFF_save_fm DFF_W1272(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25104));
DFF_save_fm DFF_W1273(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25114));
DFF_save_fm DFF_W1274(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25124));
DFF_save_fm DFF_W1275(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25204));
DFF_save_fm DFF_W1276(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25214));
DFF_save_fm DFF_W1277(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25224));
DFF_save_fm DFF_W1278(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25005));
DFF_save_fm DFF_W1279(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25015));
DFF_save_fm DFF_W1280(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25025));
DFF_save_fm DFF_W1281(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25105));
DFF_save_fm DFF_W1282(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25115));
DFF_save_fm DFF_W1283(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25125));
DFF_save_fm DFF_W1284(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25205));
DFF_save_fm DFF_W1285(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25215));
DFF_save_fm DFF_W1286(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25225));
DFF_save_fm DFF_W1287(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25006));
DFF_save_fm DFF_W1288(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25016));
DFF_save_fm DFF_W1289(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25026));
DFF_save_fm DFF_W1290(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25106));
DFF_save_fm DFF_W1291(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25116));
DFF_save_fm DFF_W1292(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25126));
DFF_save_fm DFF_W1293(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25206));
DFF_save_fm DFF_W1294(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25216));
DFF_save_fm DFF_W1295(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25226));
DFF_save_fm DFF_W1296(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25007));
DFF_save_fm DFF_W1297(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25017));
DFF_save_fm DFF_W1298(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25027));
DFF_save_fm DFF_W1299(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25107));
DFF_save_fm DFF_W1300(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25117));
DFF_save_fm DFF_W1301(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25127));
DFF_save_fm DFF_W1302(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25207));
DFF_save_fm DFF_W1303(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25217));
DFF_save_fm DFF_W1304(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25227));
DFF_save_fm DFF_W1305(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25008));
DFF_save_fm DFF_W1306(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25018));
DFF_save_fm DFF_W1307(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25028));
DFF_save_fm DFF_W1308(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25108));
DFF_save_fm DFF_W1309(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25118));
DFF_save_fm DFF_W1310(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25128));
DFF_save_fm DFF_W1311(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25208));
DFF_save_fm DFF_W1312(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25218));
DFF_save_fm DFF_W1313(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25228));
DFF_save_fm DFF_W1314(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25009));
DFF_save_fm DFF_W1315(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25019));
DFF_save_fm DFF_W1316(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25029));
DFF_save_fm DFF_W1317(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25109));
DFF_save_fm DFF_W1318(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25119));
DFF_save_fm DFF_W1319(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25129));
DFF_save_fm DFF_W1320(.clk(clk),.rstn(rstn),.reset_value(0),.q(W25209));
DFF_save_fm DFF_W1321(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25219));
DFF_save_fm DFF_W1322(.clk(clk),.rstn(rstn),.reset_value(1),.q(W25229));
DFF_save_fm DFF_W1323(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2500A));
DFF_save_fm DFF_W1324(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2501A));
DFF_save_fm DFF_W1325(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2502A));
DFF_save_fm DFF_W1326(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2510A));
DFF_save_fm DFF_W1327(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2511A));
DFF_save_fm DFF_W1328(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2512A));
DFF_save_fm DFF_W1329(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2520A));
DFF_save_fm DFF_W1330(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2521A));
DFF_save_fm DFF_W1331(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2522A));
DFF_save_fm DFF_W1332(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2500B));
DFF_save_fm DFF_W1333(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2501B));
DFF_save_fm DFF_W1334(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2502B));
DFF_save_fm DFF_W1335(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2510B));
DFF_save_fm DFF_W1336(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2511B));
DFF_save_fm DFF_W1337(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2512B));
DFF_save_fm DFF_W1338(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2520B));
DFF_save_fm DFF_W1339(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2521B));
DFF_save_fm DFF_W1340(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2522B));
DFF_save_fm DFF_W1341(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2500C));
DFF_save_fm DFF_W1342(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2501C));
DFF_save_fm DFF_W1343(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2502C));
DFF_save_fm DFF_W1344(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2510C));
DFF_save_fm DFF_W1345(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2511C));
DFF_save_fm DFF_W1346(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2512C));
DFF_save_fm DFF_W1347(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2520C));
DFF_save_fm DFF_W1348(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2521C));
DFF_save_fm DFF_W1349(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2522C));
DFF_save_fm DFF_W1350(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2500D));
DFF_save_fm DFF_W1351(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2501D));
DFF_save_fm DFF_W1352(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2502D));
DFF_save_fm DFF_W1353(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2510D));
DFF_save_fm DFF_W1354(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2511D));
DFF_save_fm DFF_W1355(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2512D));
DFF_save_fm DFF_W1356(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2520D));
DFF_save_fm DFF_W1357(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2521D));
DFF_save_fm DFF_W1358(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2522D));
DFF_save_fm DFF_W1359(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2500E));
DFF_save_fm DFF_W1360(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2501E));
DFF_save_fm DFF_W1361(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2502E));
DFF_save_fm DFF_W1362(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2510E));
DFF_save_fm DFF_W1363(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2511E));
DFF_save_fm DFF_W1364(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2512E));
DFF_save_fm DFF_W1365(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2520E));
DFF_save_fm DFF_W1366(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2521E));
DFF_save_fm DFF_W1367(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2522E));
DFF_save_fm DFF_W1368(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2500F));
DFF_save_fm DFF_W1369(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2501F));
DFF_save_fm DFF_W1370(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2502F));
DFF_save_fm DFF_W1371(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2510F));
DFF_save_fm DFF_W1372(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2511F));
DFF_save_fm DFF_W1373(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2512F));
DFF_save_fm DFF_W1374(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2520F));
DFF_save_fm DFF_W1375(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2521F));
DFF_save_fm DFF_W1376(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2522F));
DFF_save_fm DFF_W1377(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26000));
DFF_save_fm DFF_W1378(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26010));
DFF_save_fm DFF_W1379(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26020));
DFF_save_fm DFF_W1380(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26100));
DFF_save_fm DFF_W1381(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26110));
DFF_save_fm DFF_W1382(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26120));
DFF_save_fm DFF_W1383(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26200));
DFF_save_fm DFF_W1384(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26210));
DFF_save_fm DFF_W1385(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26220));
DFF_save_fm DFF_W1386(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26001));
DFF_save_fm DFF_W1387(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26011));
DFF_save_fm DFF_W1388(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26021));
DFF_save_fm DFF_W1389(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26101));
DFF_save_fm DFF_W1390(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26111));
DFF_save_fm DFF_W1391(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26121));
DFF_save_fm DFF_W1392(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26201));
DFF_save_fm DFF_W1393(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26211));
DFF_save_fm DFF_W1394(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26221));
DFF_save_fm DFF_W1395(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26002));
DFF_save_fm DFF_W1396(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26012));
DFF_save_fm DFF_W1397(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26022));
DFF_save_fm DFF_W1398(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26102));
DFF_save_fm DFF_W1399(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26112));
DFF_save_fm DFF_W1400(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26122));
DFF_save_fm DFF_W1401(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26202));
DFF_save_fm DFF_W1402(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26212));
DFF_save_fm DFF_W1403(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26222));
DFF_save_fm DFF_W1404(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26003));
DFF_save_fm DFF_W1405(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26013));
DFF_save_fm DFF_W1406(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26023));
DFF_save_fm DFF_W1407(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26103));
DFF_save_fm DFF_W1408(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26113));
DFF_save_fm DFF_W1409(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26123));
DFF_save_fm DFF_W1410(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26203));
DFF_save_fm DFF_W1411(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26213));
DFF_save_fm DFF_W1412(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26223));
DFF_save_fm DFF_W1413(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26004));
DFF_save_fm DFF_W1414(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26014));
DFF_save_fm DFF_W1415(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26024));
DFF_save_fm DFF_W1416(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26104));
DFF_save_fm DFF_W1417(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26114));
DFF_save_fm DFF_W1418(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26124));
DFF_save_fm DFF_W1419(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26204));
DFF_save_fm DFF_W1420(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26214));
DFF_save_fm DFF_W1421(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26224));
DFF_save_fm DFF_W1422(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26005));
DFF_save_fm DFF_W1423(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26015));
DFF_save_fm DFF_W1424(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26025));
DFF_save_fm DFF_W1425(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26105));
DFF_save_fm DFF_W1426(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26115));
DFF_save_fm DFF_W1427(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26125));
DFF_save_fm DFF_W1428(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26205));
DFF_save_fm DFF_W1429(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26215));
DFF_save_fm DFF_W1430(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26225));
DFF_save_fm DFF_W1431(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26006));
DFF_save_fm DFF_W1432(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26016));
DFF_save_fm DFF_W1433(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26026));
DFF_save_fm DFF_W1434(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26106));
DFF_save_fm DFF_W1435(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26116));
DFF_save_fm DFF_W1436(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26126));
DFF_save_fm DFF_W1437(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26206));
DFF_save_fm DFF_W1438(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26216));
DFF_save_fm DFF_W1439(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26226));
DFF_save_fm DFF_W1440(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26007));
DFF_save_fm DFF_W1441(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26017));
DFF_save_fm DFF_W1442(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26027));
DFF_save_fm DFF_W1443(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26107));
DFF_save_fm DFF_W1444(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26117));
DFF_save_fm DFF_W1445(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26127));
DFF_save_fm DFF_W1446(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26207));
DFF_save_fm DFF_W1447(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26217));
DFF_save_fm DFF_W1448(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26227));
DFF_save_fm DFF_W1449(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26008));
DFF_save_fm DFF_W1450(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26018));
DFF_save_fm DFF_W1451(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26028));
DFF_save_fm DFF_W1452(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26108));
DFF_save_fm DFF_W1453(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26118));
DFF_save_fm DFF_W1454(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26128));
DFF_save_fm DFF_W1455(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26208));
DFF_save_fm DFF_W1456(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26218));
DFF_save_fm DFF_W1457(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26228));
DFF_save_fm DFF_W1458(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26009));
DFF_save_fm DFF_W1459(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26019));
DFF_save_fm DFF_W1460(.clk(clk),.rstn(rstn),.reset_value(0),.q(W26029));
DFF_save_fm DFF_W1461(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26109));
DFF_save_fm DFF_W1462(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26119));
DFF_save_fm DFF_W1463(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26129));
DFF_save_fm DFF_W1464(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26209));
DFF_save_fm DFF_W1465(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26219));
DFF_save_fm DFF_W1466(.clk(clk),.rstn(rstn),.reset_value(1),.q(W26229));
DFF_save_fm DFF_W1467(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2600A));
DFF_save_fm DFF_W1468(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2601A));
DFF_save_fm DFF_W1469(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2602A));
DFF_save_fm DFF_W1470(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2610A));
DFF_save_fm DFF_W1471(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2611A));
DFF_save_fm DFF_W1472(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2612A));
DFF_save_fm DFF_W1473(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2620A));
DFF_save_fm DFF_W1474(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2621A));
DFF_save_fm DFF_W1475(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2622A));
DFF_save_fm DFF_W1476(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2600B));
DFF_save_fm DFF_W1477(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2601B));
DFF_save_fm DFF_W1478(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2602B));
DFF_save_fm DFF_W1479(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2610B));
DFF_save_fm DFF_W1480(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2611B));
DFF_save_fm DFF_W1481(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2612B));
DFF_save_fm DFF_W1482(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2620B));
DFF_save_fm DFF_W1483(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2621B));
DFF_save_fm DFF_W1484(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2622B));
DFF_save_fm DFF_W1485(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2600C));
DFF_save_fm DFF_W1486(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2601C));
DFF_save_fm DFF_W1487(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2602C));
DFF_save_fm DFF_W1488(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2610C));
DFF_save_fm DFF_W1489(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2611C));
DFF_save_fm DFF_W1490(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2612C));
DFF_save_fm DFF_W1491(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2620C));
DFF_save_fm DFF_W1492(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2621C));
DFF_save_fm DFF_W1493(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2622C));
DFF_save_fm DFF_W1494(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2600D));
DFF_save_fm DFF_W1495(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2601D));
DFF_save_fm DFF_W1496(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2602D));
DFF_save_fm DFF_W1497(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2610D));
DFF_save_fm DFF_W1498(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2611D));
DFF_save_fm DFF_W1499(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2612D));
DFF_save_fm DFF_W1500(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2620D));
DFF_save_fm DFF_W1501(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2621D));
DFF_save_fm DFF_W1502(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2622D));
DFF_save_fm DFF_W1503(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2600E));
DFF_save_fm DFF_W1504(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2601E));
DFF_save_fm DFF_W1505(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2602E));
DFF_save_fm DFF_W1506(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2610E));
DFF_save_fm DFF_W1507(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2611E));
DFF_save_fm DFF_W1508(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2612E));
DFF_save_fm DFF_W1509(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2620E));
DFF_save_fm DFF_W1510(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2621E));
DFF_save_fm DFF_W1511(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2622E));
DFF_save_fm DFF_W1512(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2600F));
DFF_save_fm DFF_W1513(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2601F));
DFF_save_fm DFF_W1514(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2602F));
DFF_save_fm DFF_W1515(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2610F));
DFF_save_fm DFF_W1516(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2611F));
DFF_save_fm DFF_W1517(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2612F));
DFF_save_fm DFF_W1518(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2620F));
DFF_save_fm DFF_W1519(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2621F));
DFF_save_fm DFF_W1520(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2622F));
DFF_save_fm DFF_W1521(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27000));
DFF_save_fm DFF_W1522(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27010));
DFF_save_fm DFF_W1523(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27020));
DFF_save_fm DFF_W1524(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27100));
DFF_save_fm DFF_W1525(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27110));
DFF_save_fm DFF_W1526(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27120));
DFF_save_fm DFF_W1527(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27200));
DFF_save_fm DFF_W1528(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27210));
DFF_save_fm DFF_W1529(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27220));
DFF_save_fm DFF_W1530(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27001));
DFF_save_fm DFF_W1531(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27011));
DFF_save_fm DFF_W1532(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27021));
DFF_save_fm DFF_W1533(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27101));
DFF_save_fm DFF_W1534(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27111));
DFF_save_fm DFF_W1535(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27121));
DFF_save_fm DFF_W1536(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27201));
DFF_save_fm DFF_W1537(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27211));
DFF_save_fm DFF_W1538(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27221));
DFF_save_fm DFF_W1539(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27002));
DFF_save_fm DFF_W1540(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27012));
DFF_save_fm DFF_W1541(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27022));
DFF_save_fm DFF_W1542(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27102));
DFF_save_fm DFF_W1543(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27112));
DFF_save_fm DFF_W1544(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27122));
DFF_save_fm DFF_W1545(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27202));
DFF_save_fm DFF_W1546(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27212));
DFF_save_fm DFF_W1547(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27222));
DFF_save_fm DFF_W1548(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27003));
DFF_save_fm DFF_W1549(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27013));
DFF_save_fm DFF_W1550(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27023));
DFF_save_fm DFF_W1551(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27103));
DFF_save_fm DFF_W1552(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27113));
DFF_save_fm DFF_W1553(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27123));
DFF_save_fm DFF_W1554(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27203));
DFF_save_fm DFF_W1555(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27213));
DFF_save_fm DFF_W1556(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27223));
DFF_save_fm DFF_W1557(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27004));
DFF_save_fm DFF_W1558(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27014));
DFF_save_fm DFF_W1559(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27024));
DFF_save_fm DFF_W1560(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27104));
DFF_save_fm DFF_W1561(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27114));
DFF_save_fm DFF_W1562(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27124));
DFF_save_fm DFF_W1563(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27204));
DFF_save_fm DFF_W1564(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27214));
DFF_save_fm DFF_W1565(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27224));
DFF_save_fm DFF_W1566(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27005));
DFF_save_fm DFF_W1567(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27015));
DFF_save_fm DFF_W1568(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27025));
DFF_save_fm DFF_W1569(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27105));
DFF_save_fm DFF_W1570(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27115));
DFF_save_fm DFF_W1571(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27125));
DFF_save_fm DFF_W1572(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27205));
DFF_save_fm DFF_W1573(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27215));
DFF_save_fm DFF_W1574(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27225));
DFF_save_fm DFF_W1575(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27006));
DFF_save_fm DFF_W1576(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27016));
DFF_save_fm DFF_W1577(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27026));
DFF_save_fm DFF_W1578(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27106));
DFF_save_fm DFF_W1579(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27116));
DFF_save_fm DFF_W1580(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27126));
DFF_save_fm DFF_W1581(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27206));
DFF_save_fm DFF_W1582(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27216));
DFF_save_fm DFF_W1583(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27226));
DFF_save_fm DFF_W1584(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27007));
DFF_save_fm DFF_W1585(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27017));
DFF_save_fm DFF_W1586(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27027));
DFF_save_fm DFF_W1587(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27107));
DFF_save_fm DFF_W1588(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27117));
DFF_save_fm DFF_W1589(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27127));
DFF_save_fm DFF_W1590(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27207));
DFF_save_fm DFF_W1591(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27217));
DFF_save_fm DFF_W1592(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27227));
DFF_save_fm DFF_W1593(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27008));
DFF_save_fm DFF_W1594(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27018));
DFF_save_fm DFF_W1595(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27028));
DFF_save_fm DFF_W1596(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27108));
DFF_save_fm DFF_W1597(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27118));
DFF_save_fm DFF_W1598(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27128));
DFF_save_fm DFF_W1599(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27208));
DFF_save_fm DFF_W1600(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27218));
DFF_save_fm DFF_W1601(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27228));
DFF_save_fm DFF_W1602(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27009));
DFF_save_fm DFF_W1603(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27019));
DFF_save_fm DFF_W1604(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27029));
DFF_save_fm DFF_W1605(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27109));
DFF_save_fm DFF_W1606(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27119));
DFF_save_fm DFF_W1607(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27129));
DFF_save_fm DFF_W1608(.clk(clk),.rstn(rstn),.reset_value(0),.q(W27209));
DFF_save_fm DFF_W1609(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27219));
DFF_save_fm DFF_W1610(.clk(clk),.rstn(rstn),.reset_value(1),.q(W27229));
DFF_save_fm DFF_W1611(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2700A));
DFF_save_fm DFF_W1612(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2701A));
DFF_save_fm DFF_W1613(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2702A));
DFF_save_fm DFF_W1614(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2710A));
DFF_save_fm DFF_W1615(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2711A));
DFF_save_fm DFF_W1616(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2712A));
DFF_save_fm DFF_W1617(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2720A));
DFF_save_fm DFF_W1618(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2721A));
DFF_save_fm DFF_W1619(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2722A));
DFF_save_fm DFF_W1620(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2700B));
DFF_save_fm DFF_W1621(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2701B));
DFF_save_fm DFF_W1622(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2702B));
DFF_save_fm DFF_W1623(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2710B));
DFF_save_fm DFF_W1624(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2711B));
DFF_save_fm DFF_W1625(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2712B));
DFF_save_fm DFF_W1626(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2720B));
DFF_save_fm DFF_W1627(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2721B));
DFF_save_fm DFF_W1628(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2722B));
DFF_save_fm DFF_W1629(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2700C));
DFF_save_fm DFF_W1630(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2701C));
DFF_save_fm DFF_W1631(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2702C));
DFF_save_fm DFF_W1632(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2710C));
DFF_save_fm DFF_W1633(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2711C));
DFF_save_fm DFF_W1634(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2712C));
DFF_save_fm DFF_W1635(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2720C));
DFF_save_fm DFF_W1636(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2721C));
DFF_save_fm DFF_W1637(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2722C));
DFF_save_fm DFF_W1638(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2700D));
DFF_save_fm DFF_W1639(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2701D));
DFF_save_fm DFF_W1640(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2702D));
DFF_save_fm DFF_W1641(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2710D));
DFF_save_fm DFF_W1642(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2711D));
DFF_save_fm DFF_W1643(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2712D));
DFF_save_fm DFF_W1644(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2720D));
DFF_save_fm DFF_W1645(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2721D));
DFF_save_fm DFF_W1646(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2722D));
DFF_save_fm DFF_W1647(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2700E));
DFF_save_fm DFF_W1648(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2701E));
DFF_save_fm DFF_W1649(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2702E));
DFF_save_fm DFF_W1650(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2710E));
DFF_save_fm DFF_W1651(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2711E));
DFF_save_fm DFF_W1652(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2712E));
DFF_save_fm DFF_W1653(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2720E));
DFF_save_fm DFF_W1654(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2721E));
DFF_save_fm DFF_W1655(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2722E));
DFF_save_fm DFF_W1656(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2700F));
DFF_save_fm DFF_W1657(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2701F));
DFF_save_fm DFF_W1658(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2702F));
DFF_save_fm DFF_W1659(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2710F));
DFF_save_fm DFF_W1660(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2711F));
DFF_save_fm DFF_W1661(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2712F));
DFF_save_fm DFF_W1662(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2720F));
DFF_save_fm DFF_W1663(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2721F));
DFF_save_fm DFF_W1664(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2722F));
DFF_save_fm DFF_W1665(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28000));
DFF_save_fm DFF_W1666(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28010));
DFF_save_fm DFF_W1667(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28020));
DFF_save_fm DFF_W1668(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28100));
DFF_save_fm DFF_W1669(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28110));
DFF_save_fm DFF_W1670(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28120));
DFF_save_fm DFF_W1671(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28200));
DFF_save_fm DFF_W1672(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28210));
DFF_save_fm DFF_W1673(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28220));
DFF_save_fm DFF_W1674(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28001));
DFF_save_fm DFF_W1675(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28011));
DFF_save_fm DFF_W1676(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28021));
DFF_save_fm DFF_W1677(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28101));
DFF_save_fm DFF_W1678(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28111));
DFF_save_fm DFF_W1679(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28121));
DFF_save_fm DFF_W1680(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28201));
DFF_save_fm DFF_W1681(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28211));
DFF_save_fm DFF_W1682(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28221));
DFF_save_fm DFF_W1683(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28002));
DFF_save_fm DFF_W1684(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28012));
DFF_save_fm DFF_W1685(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28022));
DFF_save_fm DFF_W1686(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28102));
DFF_save_fm DFF_W1687(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28112));
DFF_save_fm DFF_W1688(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28122));
DFF_save_fm DFF_W1689(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28202));
DFF_save_fm DFF_W1690(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28212));
DFF_save_fm DFF_W1691(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28222));
DFF_save_fm DFF_W1692(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28003));
DFF_save_fm DFF_W1693(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28013));
DFF_save_fm DFF_W1694(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28023));
DFF_save_fm DFF_W1695(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28103));
DFF_save_fm DFF_W1696(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28113));
DFF_save_fm DFF_W1697(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28123));
DFF_save_fm DFF_W1698(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28203));
DFF_save_fm DFF_W1699(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28213));
DFF_save_fm DFF_W1700(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28223));
DFF_save_fm DFF_W1701(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28004));
DFF_save_fm DFF_W1702(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28014));
DFF_save_fm DFF_W1703(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28024));
DFF_save_fm DFF_W1704(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28104));
DFF_save_fm DFF_W1705(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28114));
DFF_save_fm DFF_W1706(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28124));
DFF_save_fm DFF_W1707(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28204));
DFF_save_fm DFF_W1708(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28214));
DFF_save_fm DFF_W1709(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28224));
DFF_save_fm DFF_W1710(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28005));
DFF_save_fm DFF_W1711(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28015));
DFF_save_fm DFF_W1712(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28025));
DFF_save_fm DFF_W1713(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28105));
DFF_save_fm DFF_W1714(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28115));
DFF_save_fm DFF_W1715(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28125));
DFF_save_fm DFF_W1716(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28205));
DFF_save_fm DFF_W1717(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28215));
DFF_save_fm DFF_W1718(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28225));
DFF_save_fm DFF_W1719(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28006));
DFF_save_fm DFF_W1720(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28016));
DFF_save_fm DFF_W1721(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28026));
DFF_save_fm DFF_W1722(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28106));
DFF_save_fm DFF_W1723(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28116));
DFF_save_fm DFF_W1724(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28126));
DFF_save_fm DFF_W1725(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28206));
DFF_save_fm DFF_W1726(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28216));
DFF_save_fm DFF_W1727(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28226));
DFF_save_fm DFF_W1728(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28007));
DFF_save_fm DFF_W1729(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28017));
DFF_save_fm DFF_W1730(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28027));
DFF_save_fm DFF_W1731(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28107));
DFF_save_fm DFF_W1732(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28117));
DFF_save_fm DFF_W1733(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28127));
DFF_save_fm DFF_W1734(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28207));
DFF_save_fm DFF_W1735(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28217));
DFF_save_fm DFF_W1736(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28227));
DFF_save_fm DFF_W1737(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28008));
DFF_save_fm DFF_W1738(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28018));
DFF_save_fm DFF_W1739(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28028));
DFF_save_fm DFF_W1740(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28108));
DFF_save_fm DFF_W1741(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28118));
DFF_save_fm DFF_W1742(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28128));
DFF_save_fm DFF_W1743(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28208));
DFF_save_fm DFF_W1744(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28218));
DFF_save_fm DFF_W1745(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28228));
DFF_save_fm DFF_W1746(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28009));
DFF_save_fm DFF_W1747(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28019));
DFF_save_fm DFF_W1748(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28029));
DFF_save_fm DFF_W1749(.clk(clk),.rstn(rstn),.reset_value(0),.q(W28109));
DFF_save_fm DFF_W1750(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28119));
DFF_save_fm DFF_W1751(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28129));
DFF_save_fm DFF_W1752(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28209));
DFF_save_fm DFF_W1753(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28219));
DFF_save_fm DFF_W1754(.clk(clk),.rstn(rstn),.reset_value(1),.q(W28229));
DFF_save_fm DFF_W1755(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2800A));
DFF_save_fm DFF_W1756(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2801A));
DFF_save_fm DFF_W1757(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2802A));
DFF_save_fm DFF_W1758(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2810A));
DFF_save_fm DFF_W1759(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2811A));
DFF_save_fm DFF_W1760(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2812A));
DFF_save_fm DFF_W1761(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2820A));
DFF_save_fm DFF_W1762(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2821A));
DFF_save_fm DFF_W1763(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2822A));
DFF_save_fm DFF_W1764(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2800B));
DFF_save_fm DFF_W1765(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2801B));
DFF_save_fm DFF_W1766(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2802B));
DFF_save_fm DFF_W1767(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2810B));
DFF_save_fm DFF_W1768(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2811B));
DFF_save_fm DFF_W1769(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2812B));
DFF_save_fm DFF_W1770(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2820B));
DFF_save_fm DFF_W1771(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2821B));
DFF_save_fm DFF_W1772(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2822B));
DFF_save_fm DFF_W1773(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2800C));
DFF_save_fm DFF_W1774(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2801C));
DFF_save_fm DFF_W1775(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2802C));
DFF_save_fm DFF_W1776(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2810C));
DFF_save_fm DFF_W1777(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2811C));
DFF_save_fm DFF_W1778(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2812C));
DFF_save_fm DFF_W1779(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2820C));
DFF_save_fm DFF_W1780(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2821C));
DFF_save_fm DFF_W1781(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2822C));
DFF_save_fm DFF_W1782(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2800D));
DFF_save_fm DFF_W1783(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2801D));
DFF_save_fm DFF_W1784(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2802D));
DFF_save_fm DFF_W1785(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2810D));
DFF_save_fm DFF_W1786(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2811D));
DFF_save_fm DFF_W1787(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2812D));
DFF_save_fm DFF_W1788(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2820D));
DFF_save_fm DFF_W1789(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2821D));
DFF_save_fm DFF_W1790(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2822D));
DFF_save_fm DFF_W1791(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2800E));
DFF_save_fm DFF_W1792(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2801E));
DFF_save_fm DFF_W1793(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2802E));
DFF_save_fm DFF_W1794(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2810E));
DFF_save_fm DFF_W1795(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2811E));
DFF_save_fm DFF_W1796(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2812E));
DFF_save_fm DFF_W1797(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2820E));
DFF_save_fm DFF_W1798(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2821E));
DFF_save_fm DFF_W1799(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2822E));
DFF_save_fm DFF_W1800(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2800F));
DFF_save_fm DFF_W1801(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2801F));
DFF_save_fm DFF_W1802(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2802F));
DFF_save_fm DFF_W1803(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2810F));
DFF_save_fm DFF_W1804(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2811F));
DFF_save_fm DFF_W1805(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2812F));
DFF_save_fm DFF_W1806(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2820F));
DFF_save_fm DFF_W1807(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2821F));
DFF_save_fm DFF_W1808(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2822F));
DFF_save_fm DFF_W1809(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29000));
DFF_save_fm DFF_W1810(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29010));
DFF_save_fm DFF_W1811(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29020));
DFF_save_fm DFF_W1812(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29100));
DFF_save_fm DFF_W1813(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29110));
DFF_save_fm DFF_W1814(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29120));
DFF_save_fm DFF_W1815(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29200));
DFF_save_fm DFF_W1816(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29210));
DFF_save_fm DFF_W1817(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29220));
DFF_save_fm DFF_W1818(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29001));
DFF_save_fm DFF_W1819(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29011));
DFF_save_fm DFF_W1820(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29021));
DFF_save_fm DFF_W1821(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29101));
DFF_save_fm DFF_W1822(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29111));
DFF_save_fm DFF_W1823(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29121));
DFF_save_fm DFF_W1824(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29201));
DFF_save_fm DFF_W1825(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29211));
DFF_save_fm DFF_W1826(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29221));
DFF_save_fm DFF_W1827(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29002));
DFF_save_fm DFF_W1828(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29012));
DFF_save_fm DFF_W1829(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29022));
DFF_save_fm DFF_W1830(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29102));
DFF_save_fm DFF_W1831(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29112));
DFF_save_fm DFF_W1832(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29122));
DFF_save_fm DFF_W1833(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29202));
DFF_save_fm DFF_W1834(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29212));
DFF_save_fm DFF_W1835(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29222));
DFF_save_fm DFF_W1836(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29003));
DFF_save_fm DFF_W1837(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29013));
DFF_save_fm DFF_W1838(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29023));
DFF_save_fm DFF_W1839(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29103));
DFF_save_fm DFF_W1840(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29113));
DFF_save_fm DFF_W1841(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29123));
DFF_save_fm DFF_W1842(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29203));
DFF_save_fm DFF_W1843(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29213));
DFF_save_fm DFF_W1844(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29223));
DFF_save_fm DFF_W1845(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29004));
DFF_save_fm DFF_W1846(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29014));
DFF_save_fm DFF_W1847(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29024));
DFF_save_fm DFF_W1848(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29104));
DFF_save_fm DFF_W1849(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29114));
DFF_save_fm DFF_W1850(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29124));
DFF_save_fm DFF_W1851(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29204));
DFF_save_fm DFF_W1852(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29214));
DFF_save_fm DFF_W1853(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29224));
DFF_save_fm DFF_W1854(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29005));
DFF_save_fm DFF_W1855(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29015));
DFF_save_fm DFF_W1856(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29025));
DFF_save_fm DFF_W1857(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29105));
DFF_save_fm DFF_W1858(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29115));
DFF_save_fm DFF_W1859(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29125));
DFF_save_fm DFF_W1860(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29205));
DFF_save_fm DFF_W1861(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29215));
DFF_save_fm DFF_W1862(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29225));
DFF_save_fm DFF_W1863(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29006));
DFF_save_fm DFF_W1864(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29016));
DFF_save_fm DFF_W1865(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29026));
DFF_save_fm DFF_W1866(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29106));
DFF_save_fm DFF_W1867(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29116));
DFF_save_fm DFF_W1868(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29126));
DFF_save_fm DFF_W1869(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29206));
DFF_save_fm DFF_W1870(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29216));
DFF_save_fm DFF_W1871(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29226));
DFF_save_fm DFF_W1872(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29007));
DFF_save_fm DFF_W1873(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29017));
DFF_save_fm DFF_W1874(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29027));
DFF_save_fm DFF_W1875(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29107));
DFF_save_fm DFF_W1876(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29117));
DFF_save_fm DFF_W1877(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29127));
DFF_save_fm DFF_W1878(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29207));
DFF_save_fm DFF_W1879(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29217));
DFF_save_fm DFF_W1880(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29227));
DFF_save_fm DFF_W1881(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29008));
DFF_save_fm DFF_W1882(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29018));
DFF_save_fm DFF_W1883(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29028));
DFF_save_fm DFF_W1884(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29108));
DFF_save_fm DFF_W1885(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29118));
DFF_save_fm DFF_W1886(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29128));
DFF_save_fm DFF_W1887(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29208));
DFF_save_fm DFF_W1888(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29218));
DFF_save_fm DFF_W1889(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29228));
DFF_save_fm DFF_W1890(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29009));
DFF_save_fm DFF_W1891(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29019));
DFF_save_fm DFF_W1892(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29029));
DFF_save_fm DFF_W1893(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29109));
DFF_save_fm DFF_W1894(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29119));
DFF_save_fm DFF_W1895(.clk(clk),.rstn(rstn),.reset_value(1),.q(W29129));
DFF_save_fm DFF_W1896(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29209));
DFF_save_fm DFF_W1897(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29219));
DFF_save_fm DFF_W1898(.clk(clk),.rstn(rstn),.reset_value(0),.q(W29229));
DFF_save_fm DFF_W1899(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2900A));
DFF_save_fm DFF_W1900(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2901A));
DFF_save_fm DFF_W1901(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2902A));
DFF_save_fm DFF_W1902(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2910A));
DFF_save_fm DFF_W1903(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2911A));
DFF_save_fm DFF_W1904(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2912A));
DFF_save_fm DFF_W1905(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2920A));
DFF_save_fm DFF_W1906(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2921A));
DFF_save_fm DFF_W1907(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2922A));
DFF_save_fm DFF_W1908(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2900B));
DFF_save_fm DFF_W1909(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2901B));
DFF_save_fm DFF_W1910(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2902B));
DFF_save_fm DFF_W1911(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2910B));
DFF_save_fm DFF_W1912(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2911B));
DFF_save_fm DFF_W1913(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2912B));
DFF_save_fm DFF_W1914(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2920B));
DFF_save_fm DFF_W1915(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2921B));
DFF_save_fm DFF_W1916(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2922B));
DFF_save_fm DFF_W1917(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2900C));
DFF_save_fm DFF_W1918(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2901C));
DFF_save_fm DFF_W1919(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2902C));
DFF_save_fm DFF_W1920(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2910C));
DFF_save_fm DFF_W1921(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2911C));
DFF_save_fm DFF_W1922(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2912C));
DFF_save_fm DFF_W1923(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2920C));
DFF_save_fm DFF_W1924(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2921C));
DFF_save_fm DFF_W1925(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2922C));
DFF_save_fm DFF_W1926(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2900D));
DFF_save_fm DFF_W1927(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2901D));
DFF_save_fm DFF_W1928(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2902D));
DFF_save_fm DFF_W1929(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2910D));
DFF_save_fm DFF_W1930(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2911D));
DFF_save_fm DFF_W1931(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2912D));
DFF_save_fm DFF_W1932(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2920D));
DFF_save_fm DFF_W1933(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2921D));
DFF_save_fm DFF_W1934(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2922D));
DFF_save_fm DFF_W1935(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2900E));
DFF_save_fm DFF_W1936(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2901E));
DFF_save_fm DFF_W1937(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2902E));
DFF_save_fm DFF_W1938(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2910E));
DFF_save_fm DFF_W1939(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2911E));
DFF_save_fm DFF_W1940(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2912E));
DFF_save_fm DFF_W1941(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2920E));
DFF_save_fm DFF_W1942(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2921E));
DFF_save_fm DFF_W1943(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2922E));
DFF_save_fm DFF_W1944(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2900F));
DFF_save_fm DFF_W1945(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2901F));
DFF_save_fm DFF_W1946(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2902F));
DFF_save_fm DFF_W1947(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2910F));
DFF_save_fm DFF_W1948(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2911F));
DFF_save_fm DFF_W1949(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2912F));
DFF_save_fm DFF_W1950(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2920F));
DFF_save_fm DFF_W1951(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2921F));
DFF_save_fm DFF_W1952(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2922F));
DFF_save_fm DFF_W1953(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A000));
DFF_save_fm DFF_W1954(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A010));
DFF_save_fm DFF_W1955(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A020));
DFF_save_fm DFF_W1956(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A100));
DFF_save_fm DFF_W1957(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A110));
DFF_save_fm DFF_W1958(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A120));
DFF_save_fm DFF_W1959(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A200));
DFF_save_fm DFF_W1960(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A210));
DFF_save_fm DFF_W1961(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A220));
DFF_save_fm DFF_W1962(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A001));
DFF_save_fm DFF_W1963(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A011));
DFF_save_fm DFF_W1964(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A021));
DFF_save_fm DFF_W1965(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A101));
DFF_save_fm DFF_W1966(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A111));
DFF_save_fm DFF_W1967(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A121));
DFF_save_fm DFF_W1968(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A201));
DFF_save_fm DFF_W1969(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A211));
DFF_save_fm DFF_W1970(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A221));
DFF_save_fm DFF_W1971(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A002));
DFF_save_fm DFF_W1972(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A012));
DFF_save_fm DFF_W1973(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A022));
DFF_save_fm DFF_W1974(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A102));
DFF_save_fm DFF_W1975(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A112));
DFF_save_fm DFF_W1976(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A122));
DFF_save_fm DFF_W1977(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A202));
DFF_save_fm DFF_W1978(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A212));
DFF_save_fm DFF_W1979(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A222));
DFF_save_fm DFF_W1980(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A003));
DFF_save_fm DFF_W1981(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A013));
DFF_save_fm DFF_W1982(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A023));
DFF_save_fm DFF_W1983(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A103));
DFF_save_fm DFF_W1984(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A113));
DFF_save_fm DFF_W1985(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A123));
DFF_save_fm DFF_W1986(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A203));
DFF_save_fm DFF_W1987(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A213));
DFF_save_fm DFF_W1988(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A223));
DFF_save_fm DFF_W1989(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A004));
DFF_save_fm DFF_W1990(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A014));
DFF_save_fm DFF_W1991(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A024));
DFF_save_fm DFF_W1992(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A104));
DFF_save_fm DFF_W1993(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A114));
DFF_save_fm DFF_W1994(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A124));
DFF_save_fm DFF_W1995(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A204));
DFF_save_fm DFF_W1996(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A214));
DFF_save_fm DFF_W1997(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A224));
DFF_save_fm DFF_W1998(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A005));
DFF_save_fm DFF_W1999(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A015));
DFF_save_fm DFF_W2000(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A025));
DFF_save_fm DFF_W2001(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A105));
DFF_save_fm DFF_W2002(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A115));
DFF_save_fm DFF_W2003(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A125));
DFF_save_fm DFF_W2004(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A205));
DFF_save_fm DFF_W2005(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A215));
DFF_save_fm DFF_W2006(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A225));
DFF_save_fm DFF_W2007(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A006));
DFF_save_fm DFF_W2008(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A016));
DFF_save_fm DFF_W2009(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A026));
DFF_save_fm DFF_W2010(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A106));
DFF_save_fm DFF_W2011(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A116));
DFF_save_fm DFF_W2012(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A126));
DFF_save_fm DFF_W2013(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A206));
DFF_save_fm DFF_W2014(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A216));
DFF_save_fm DFF_W2015(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A226));
DFF_save_fm DFF_W2016(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A007));
DFF_save_fm DFF_W2017(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A017));
DFF_save_fm DFF_W2018(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A027));
DFF_save_fm DFF_W2019(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A107));
DFF_save_fm DFF_W2020(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A117));
DFF_save_fm DFF_W2021(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A127));
DFF_save_fm DFF_W2022(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A207));
DFF_save_fm DFF_W2023(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A217));
DFF_save_fm DFF_W2024(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A227));
DFF_save_fm DFF_W2025(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A008));
DFF_save_fm DFF_W2026(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A018));
DFF_save_fm DFF_W2027(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A028));
DFF_save_fm DFF_W2028(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A108));
DFF_save_fm DFF_W2029(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A118));
DFF_save_fm DFF_W2030(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A128));
DFF_save_fm DFF_W2031(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A208));
DFF_save_fm DFF_W2032(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A218));
DFF_save_fm DFF_W2033(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A228));
DFF_save_fm DFF_W2034(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A009));
DFF_save_fm DFF_W2035(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A019));
DFF_save_fm DFF_W2036(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A029));
DFF_save_fm DFF_W2037(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A109));
DFF_save_fm DFF_W2038(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A119));
DFF_save_fm DFF_W2039(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A129));
DFF_save_fm DFF_W2040(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A209));
DFF_save_fm DFF_W2041(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A219));
DFF_save_fm DFF_W2042(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A229));
DFF_save_fm DFF_W2043(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A00A));
DFF_save_fm DFF_W2044(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A01A));
DFF_save_fm DFF_W2045(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A02A));
DFF_save_fm DFF_W2046(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A10A));
DFF_save_fm DFF_W2047(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A11A));
DFF_save_fm DFF_W2048(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A12A));
DFF_save_fm DFF_W2049(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A20A));
DFF_save_fm DFF_W2050(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A21A));
DFF_save_fm DFF_W2051(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A22A));
DFF_save_fm DFF_W2052(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A00B));
DFF_save_fm DFF_W2053(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A01B));
DFF_save_fm DFF_W2054(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A02B));
DFF_save_fm DFF_W2055(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A10B));
DFF_save_fm DFF_W2056(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A11B));
DFF_save_fm DFF_W2057(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A12B));
DFF_save_fm DFF_W2058(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A20B));
DFF_save_fm DFF_W2059(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A21B));
DFF_save_fm DFF_W2060(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A22B));
DFF_save_fm DFF_W2061(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A00C));
DFF_save_fm DFF_W2062(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A01C));
DFF_save_fm DFF_W2063(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A02C));
DFF_save_fm DFF_W2064(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A10C));
DFF_save_fm DFF_W2065(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A11C));
DFF_save_fm DFF_W2066(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A12C));
DFF_save_fm DFF_W2067(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A20C));
DFF_save_fm DFF_W2068(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A21C));
DFF_save_fm DFF_W2069(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A22C));
DFF_save_fm DFF_W2070(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A00D));
DFF_save_fm DFF_W2071(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A01D));
DFF_save_fm DFF_W2072(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A02D));
DFF_save_fm DFF_W2073(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A10D));
DFF_save_fm DFF_W2074(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A11D));
DFF_save_fm DFF_W2075(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A12D));
DFF_save_fm DFF_W2076(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A20D));
DFF_save_fm DFF_W2077(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A21D));
DFF_save_fm DFF_W2078(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A22D));
DFF_save_fm DFF_W2079(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A00E));
DFF_save_fm DFF_W2080(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A01E));
DFF_save_fm DFF_W2081(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A02E));
DFF_save_fm DFF_W2082(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A10E));
DFF_save_fm DFF_W2083(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A11E));
DFF_save_fm DFF_W2084(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A12E));
DFF_save_fm DFF_W2085(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A20E));
DFF_save_fm DFF_W2086(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A21E));
DFF_save_fm DFF_W2087(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A22E));
DFF_save_fm DFF_W2088(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A00F));
DFF_save_fm DFF_W2089(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A01F));
DFF_save_fm DFF_W2090(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A02F));
DFF_save_fm DFF_W2091(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A10F));
DFF_save_fm DFF_W2092(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A11F));
DFF_save_fm DFF_W2093(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A12F));
DFF_save_fm DFF_W2094(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A20F));
DFF_save_fm DFF_W2095(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2A21F));
DFF_save_fm DFF_W2096(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2A22F));
DFF_save_fm DFF_W2097(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B000));
DFF_save_fm DFF_W2098(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B010));
DFF_save_fm DFF_W2099(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B020));
DFF_save_fm DFF_W2100(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B100));
DFF_save_fm DFF_W2101(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B110));
DFF_save_fm DFF_W2102(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B120));
DFF_save_fm DFF_W2103(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B200));
DFF_save_fm DFF_W2104(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B210));
DFF_save_fm DFF_W2105(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B220));
DFF_save_fm DFF_W2106(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B001));
DFF_save_fm DFF_W2107(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B011));
DFF_save_fm DFF_W2108(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B021));
DFF_save_fm DFF_W2109(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B101));
DFF_save_fm DFF_W2110(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B111));
DFF_save_fm DFF_W2111(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B121));
DFF_save_fm DFF_W2112(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B201));
DFF_save_fm DFF_W2113(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B211));
DFF_save_fm DFF_W2114(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B221));
DFF_save_fm DFF_W2115(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B002));
DFF_save_fm DFF_W2116(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B012));
DFF_save_fm DFF_W2117(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B022));
DFF_save_fm DFF_W2118(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B102));
DFF_save_fm DFF_W2119(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B112));
DFF_save_fm DFF_W2120(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B122));
DFF_save_fm DFF_W2121(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B202));
DFF_save_fm DFF_W2122(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B212));
DFF_save_fm DFF_W2123(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B222));
DFF_save_fm DFF_W2124(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B003));
DFF_save_fm DFF_W2125(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B013));
DFF_save_fm DFF_W2126(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B023));
DFF_save_fm DFF_W2127(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B103));
DFF_save_fm DFF_W2128(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B113));
DFF_save_fm DFF_W2129(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B123));
DFF_save_fm DFF_W2130(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B203));
DFF_save_fm DFF_W2131(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B213));
DFF_save_fm DFF_W2132(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B223));
DFF_save_fm DFF_W2133(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B004));
DFF_save_fm DFF_W2134(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B014));
DFF_save_fm DFF_W2135(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B024));
DFF_save_fm DFF_W2136(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B104));
DFF_save_fm DFF_W2137(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B114));
DFF_save_fm DFF_W2138(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B124));
DFF_save_fm DFF_W2139(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B204));
DFF_save_fm DFF_W2140(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B214));
DFF_save_fm DFF_W2141(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B224));
DFF_save_fm DFF_W2142(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B005));
DFF_save_fm DFF_W2143(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B015));
DFF_save_fm DFF_W2144(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B025));
DFF_save_fm DFF_W2145(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B105));
DFF_save_fm DFF_W2146(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B115));
DFF_save_fm DFF_W2147(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B125));
DFF_save_fm DFF_W2148(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B205));
DFF_save_fm DFF_W2149(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B215));
DFF_save_fm DFF_W2150(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B225));
DFF_save_fm DFF_W2151(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B006));
DFF_save_fm DFF_W2152(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B016));
DFF_save_fm DFF_W2153(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B026));
DFF_save_fm DFF_W2154(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B106));
DFF_save_fm DFF_W2155(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B116));
DFF_save_fm DFF_W2156(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B126));
DFF_save_fm DFF_W2157(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B206));
DFF_save_fm DFF_W2158(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B216));
DFF_save_fm DFF_W2159(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B226));
DFF_save_fm DFF_W2160(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B007));
DFF_save_fm DFF_W2161(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B017));
DFF_save_fm DFF_W2162(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B027));
DFF_save_fm DFF_W2163(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B107));
DFF_save_fm DFF_W2164(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B117));
DFF_save_fm DFF_W2165(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B127));
DFF_save_fm DFF_W2166(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B207));
DFF_save_fm DFF_W2167(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B217));
DFF_save_fm DFF_W2168(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B227));
DFF_save_fm DFF_W2169(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B008));
DFF_save_fm DFF_W2170(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B018));
DFF_save_fm DFF_W2171(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B028));
DFF_save_fm DFF_W2172(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B108));
DFF_save_fm DFF_W2173(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B118));
DFF_save_fm DFF_W2174(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B128));
DFF_save_fm DFF_W2175(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B208));
DFF_save_fm DFF_W2176(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B218));
DFF_save_fm DFF_W2177(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B228));
DFF_save_fm DFF_W2178(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B009));
DFF_save_fm DFF_W2179(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B019));
DFF_save_fm DFF_W2180(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B029));
DFF_save_fm DFF_W2181(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B109));
DFF_save_fm DFF_W2182(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B119));
DFF_save_fm DFF_W2183(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B129));
DFF_save_fm DFF_W2184(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B209));
DFF_save_fm DFF_W2185(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B219));
DFF_save_fm DFF_W2186(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B229));
DFF_save_fm DFF_W2187(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B00A));
DFF_save_fm DFF_W2188(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B01A));
DFF_save_fm DFF_W2189(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B02A));
DFF_save_fm DFF_W2190(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B10A));
DFF_save_fm DFF_W2191(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B11A));
DFF_save_fm DFF_W2192(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B12A));
DFF_save_fm DFF_W2193(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B20A));
DFF_save_fm DFF_W2194(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B21A));
DFF_save_fm DFF_W2195(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B22A));
DFF_save_fm DFF_W2196(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B00B));
DFF_save_fm DFF_W2197(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B01B));
DFF_save_fm DFF_W2198(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B02B));
DFF_save_fm DFF_W2199(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B10B));
DFF_save_fm DFF_W2200(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B11B));
DFF_save_fm DFF_W2201(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B12B));
DFF_save_fm DFF_W2202(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B20B));
DFF_save_fm DFF_W2203(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B21B));
DFF_save_fm DFF_W2204(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B22B));
DFF_save_fm DFF_W2205(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B00C));
DFF_save_fm DFF_W2206(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B01C));
DFF_save_fm DFF_W2207(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B02C));
DFF_save_fm DFF_W2208(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B10C));
DFF_save_fm DFF_W2209(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B11C));
DFF_save_fm DFF_W2210(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B12C));
DFF_save_fm DFF_W2211(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B20C));
DFF_save_fm DFF_W2212(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B21C));
DFF_save_fm DFF_W2213(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B22C));
DFF_save_fm DFF_W2214(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B00D));
DFF_save_fm DFF_W2215(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B01D));
DFF_save_fm DFF_W2216(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B02D));
DFF_save_fm DFF_W2217(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B10D));
DFF_save_fm DFF_W2218(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B11D));
DFF_save_fm DFF_W2219(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B12D));
DFF_save_fm DFF_W2220(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B20D));
DFF_save_fm DFF_W2221(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B21D));
DFF_save_fm DFF_W2222(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B22D));
DFF_save_fm DFF_W2223(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B00E));
DFF_save_fm DFF_W2224(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B01E));
DFF_save_fm DFF_W2225(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B02E));
DFF_save_fm DFF_W2226(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B10E));
DFF_save_fm DFF_W2227(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B11E));
DFF_save_fm DFF_W2228(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B12E));
DFF_save_fm DFF_W2229(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B20E));
DFF_save_fm DFF_W2230(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B21E));
DFF_save_fm DFF_W2231(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B22E));
DFF_save_fm DFF_W2232(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B00F));
DFF_save_fm DFF_W2233(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B01F));
DFF_save_fm DFF_W2234(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B02F));
DFF_save_fm DFF_W2235(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B10F));
DFF_save_fm DFF_W2236(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B11F));
DFF_save_fm DFF_W2237(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B12F));
DFF_save_fm DFF_W2238(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2B20F));
DFF_save_fm DFF_W2239(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B21F));
DFF_save_fm DFF_W2240(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2B22F));
DFF_save_fm DFF_W2241(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C000));
DFF_save_fm DFF_W2242(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C010));
DFF_save_fm DFF_W2243(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C020));
DFF_save_fm DFF_W2244(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C100));
DFF_save_fm DFF_W2245(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C110));
DFF_save_fm DFF_W2246(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C120));
DFF_save_fm DFF_W2247(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C200));
DFF_save_fm DFF_W2248(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C210));
DFF_save_fm DFF_W2249(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C220));
DFF_save_fm DFF_W2250(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C001));
DFF_save_fm DFF_W2251(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C011));
DFF_save_fm DFF_W2252(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C021));
DFF_save_fm DFF_W2253(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C101));
DFF_save_fm DFF_W2254(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C111));
DFF_save_fm DFF_W2255(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C121));
DFF_save_fm DFF_W2256(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C201));
DFF_save_fm DFF_W2257(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C211));
DFF_save_fm DFF_W2258(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C221));
DFF_save_fm DFF_W2259(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C002));
DFF_save_fm DFF_W2260(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C012));
DFF_save_fm DFF_W2261(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C022));
DFF_save_fm DFF_W2262(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C102));
DFF_save_fm DFF_W2263(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C112));
DFF_save_fm DFF_W2264(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C122));
DFF_save_fm DFF_W2265(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C202));
DFF_save_fm DFF_W2266(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C212));
DFF_save_fm DFF_W2267(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C222));
DFF_save_fm DFF_W2268(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C003));
DFF_save_fm DFF_W2269(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C013));
DFF_save_fm DFF_W2270(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C023));
DFF_save_fm DFF_W2271(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C103));
DFF_save_fm DFF_W2272(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C113));
DFF_save_fm DFF_W2273(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C123));
DFF_save_fm DFF_W2274(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C203));
DFF_save_fm DFF_W2275(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C213));
DFF_save_fm DFF_W2276(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C223));
DFF_save_fm DFF_W2277(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C004));
DFF_save_fm DFF_W2278(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C014));
DFF_save_fm DFF_W2279(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C024));
DFF_save_fm DFF_W2280(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C104));
DFF_save_fm DFF_W2281(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C114));
DFF_save_fm DFF_W2282(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C124));
DFF_save_fm DFF_W2283(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C204));
DFF_save_fm DFF_W2284(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C214));
DFF_save_fm DFF_W2285(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C224));
DFF_save_fm DFF_W2286(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C005));
DFF_save_fm DFF_W2287(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C015));
DFF_save_fm DFF_W2288(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C025));
DFF_save_fm DFF_W2289(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C105));
DFF_save_fm DFF_W2290(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C115));
DFF_save_fm DFF_W2291(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C125));
DFF_save_fm DFF_W2292(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C205));
DFF_save_fm DFF_W2293(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C215));
DFF_save_fm DFF_W2294(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C225));
DFF_save_fm DFF_W2295(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C006));
DFF_save_fm DFF_W2296(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C016));
DFF_save_fm DFF_W2297(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C026));
DFF_save_fm DFF_W2298(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C106));
DFF_save_fm DFF_W2299(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C116));
DFF_save_fm DFF_W2300(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C126));
DFF_save_fm DFF_W2301(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C206));
DFF_save_fm DFF_W2302(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C216));
DFF_save_fm DFF_W2303(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C226));
DFF_save_fm DFF_W2304(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C007));
DFF_save_fm DFF_W2305(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C017));
DFF_save_fm DFF_W2306(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C027));
DFF_save_fm DFF_W2307(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C107));
DFF_save_fm DFF_W2308(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C117));
DFF_save_fm DFF_W2309(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C127));
DFF_save_fm DFF_W2310(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C207));
DFF_save_fm DFF_W2311(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C217));
DFF_save_fm DFF_W2312(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C227));
DFF_save_fm DFF_W2313(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C008));
DFF_save_fm DFF_W2314(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C018));
DFF_save_fm DFF_W2315(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C028));
DFF_save_fm DFF_W2316(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C108));
DFF_save_fm DFF_W2317(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C118));
DFF_save_fm DFF_W2318(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C128));
DFF_save_fm DFF_W2319(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C208));
DFF_save_fm DFF_W2320(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C218));
DFF_save_fm DFF_W2321(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C228));
DFF_save_fm DFF_W2322(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C009));
DFF_save_fm DFF_W2323(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C019));
DFF_save_fm DFF_W2324(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C029));
DFF_save_fm DFF_W2325(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C109));
DFF_save_fm DFF_W2326(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C119));
DFF_save_fm DFF_W2327(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C129));
DFF_save_fm DFF_W2328(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C209));
DFF_save_fm DFF_W2329(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C219));
DFF_save_fm DFF_W2330(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C229));
DFF_save_fm DFF_W2331(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C00A));
DFF_save_fm DFF_W2332(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C01A));
DFF_save_fm DFF_W2333(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C02A));
DFF_save_fm DFF_W2334(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C10A));
DFF_save_fm DFF_W2335(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C11A));
DFF_save_fm DFF_W2336(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C12A));
DFF_save_fm DFF_W2337(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C20A));
DFF_save_fm DFF_W2338(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C21A));
DFF_save_fm DFF_W2339(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C22A));
DFF_save_fm DFF_W2340(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C00B));
DFF_save_fm DFF_W2341(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C01B));
DFF_save_fm DFF_W2342(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C02B));
DFF_save_fm DFF_W2343(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C10B));
DFF_save_fm DFF_W2344(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C11B));
DFF_save_fm DFF_W2345(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C12B));
DFF_save_fm DFF_W2346(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C20B));
DFF_save_fm DFF_W2347(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C21B));
DFF_save_fm DFF_W2348(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C22B));
DFF_save_fm DFF_W2349(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C00C));
DFF_save_fm DFF_W2350(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C01C));
DFF_save_fm DFF_W2351(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C02C));
DFF_save_fm DFF_W2352(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C10C));
DFF_save_fm DFF_W2353(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C11C));
DFF_save_fm DFF_W2354(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C12C));
DFF_save_fm DFF_W2355(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C20C));
DFF_save_fm DFF_W2356(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C21C));
DFF_save_fm DFF_W2357(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C22C));
DFF_save_fm DFF_W2358(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C00D));
DFF_save_fm DFF_W2359(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C01D));
DFF_save_fm DFF_W2360(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C02D));
DFF_save_fm DFF_W2361(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C10D));
DFF_save_fm DFF_W2362(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C11D));
DFF_save_fm DFF_W2363(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C12D));
DFF_save_fm DFF_W2364(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C20D));
DFF_save_fm DFF_W2365(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C21D));
DFF_save_fm DFF_W2366(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C22D));
DFF_save_fm DFF_W2367(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C00E));
DFF_save_fm DFF_W2368(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C01E));
DFF_save_fm DFF_W2369(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C02E));
DFF_save_fm DFF_W2370(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C10E));
DFF_save_fm DFF_W2371(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C11E));
DFF_save_fm DFF_W2372(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C12E));
DFF_save_fm DFF_W2373(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C20E));
DFF_save_fm DFF_W2374(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C21E));
DFF_save_fm DFF_W2375(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C22E));
DFF_save_fm DFF_W2376(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C00F));
DFF_save_fm DFF_W2377(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C01F));
DFF_save_fm DFF_W2378(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C02F));
DFF_save_fm DFF_W2379(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C10F));
DFF_save_fm DFF_W2380(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C11F));
DFF_save_fm DFF_W2381(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2C12F));
DFF_save_fm DFF_W2382(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C20F));
DFF_save_fm DFF_W2383(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C21F));
DFF_save_fm DFF_W2384(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2C22F));
DFF_save_fm DFF_W2385(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D000));
DFF_save_fm DFF_W2386(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D010));
DFF_save_fm DFF_W2387(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D020));
DFF_save_fm DFF_W2388(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D100));
DFF_save_fm DFF_W2389(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D110));
DFF_save_fm DFF_W2390(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D120));
DFF_save_fm DFF_W2391(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D200));
DFF_save_fm DFF_W2392(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D210));
DFF_save_fm DFF_W2393(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D220));
DFF_save_fm DFF_W2394(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D001));
DFF_save_fm DFF_W2395(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D011));
DFF_save_fm DFF_W2396(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D021));
DFF_save_fm DFF_W2397(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D101));
DFF_save_fm DFF_W2398(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D111));
DFF_save_fm DFF_W2399(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D121));
DFF_save_fm DFF_W2400(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D201));
DFF_save_fm DFF_W2401(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D211));
DFF_save_fm DFF_W2402(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D221));
DFF_save_fm DFF_W2403(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D002));
DFF_save_fm DFF_W2404(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D012));
DFF_save_fm DFF_W2405(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D022));
DFF_save_fm DFF_W2406(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D102));
DFF_save_fm DFF_W2407(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D112));
DFF_save_fm DFF_W2408(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D122));
DFF_save_fm DFF_W2409(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D202));
DFF_save_fm DFF_W2410(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D212));
DFF_save_fm DFF_W2411(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D222));
DFF_save_fm DFF_W2412(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D003));
DFF_save_fm DFF_W2413(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D013));
DFF_save_fm DFF_W2414(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D023));
DFF_save_fm DFF_W2415(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D103));
DFF_save_fm DFF_W2416(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D113));
DFF_save_fm DFF_W2417(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D123));
DFF_save_fm DFF_W2418(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D203));
DFF_save_fm DFF_W2419(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D213));
DFF_save_fm DFF_W2420(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D223));
DFF_save_fm DFF_W2421(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D004));
DFF_save_fm DFF_W2422(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D014));
DFF_save_fm DFF_W2423(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D024));
DFF_save_fm DFF_W2424(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D104));
DFF_save_fm DFF_W2425(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D114));
DFF_save_fm DFF_W2426(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D124));
DFF_save_fm DFF_W2427(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D204));
DFF_save_fm DFF_W2428(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D214));
DFF_save_fm DFF_W2429(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D224));
DFF_save_fm DFF_W2430(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D005));
DFF_save_fm DFF_W2431(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D015));
DFF_save_fm DFF_W2432(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D025));
DFF_save_fm DFF_W2433(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D105));
DFF_save_fm DFF_W2434(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D115));
DFF_save_fm DFF_W2435(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D125));
DFF_save_fm DFF_W2436(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D205));
DFF_save_fm DFF_W2437(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D215));
DFF_save_fm DFF_W2438(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D225));
DFF_save_fm DFF_W2439(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D006));
DFF_save_fm DFF_W2440(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D016));
DFF_save_fm DFF_W2441(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D026));
DFF_save_fm DFF_W2442(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D106));
DFF_save_fm DFF_W2443(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D116));
DFF_save_fm DFF_W2444(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D126));
DFF_save_fm DFF_W2445(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D206));
DFF_save_fm DFF_W2446(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D216));
DFF_save_fm DFF_W2447(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D226));
DFF_save_fm DFF_W2448(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D007));
DFF_save_fm DFF_W2449(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D017));
DFF_save_fm DFF_W2450(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D027));
DFF_save_fm DFF_W2451(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D107));
DFF_save_fm DFF_W2452(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D117));
DFF_save_fm DFF_W2453(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D127));
DFF_save_fm DFF_W2454(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D207));
DFF_save_fm DFF_W2455(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D217));
DFF_save_fm DFF_W2456(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D227));
DFF_save_fm DFF_W2457(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D008));
DFF_save_fm DFF_W2458(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D018));
DFF_save_fm DFF_W2459(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D028));
DFF_save_fm DFF_W2460(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D108));
DFF_save_fm DFF_W2461(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D118));
DFF_save_fm DFF_W2462(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D128));
DFF_save_fm DFF_W2463(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D208));
DFF_save_fm DFF_W2464(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D218));
DFF_save_fm DFF_W2465(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D228));
DFF_save_fm DFF_W2466(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D009));
DFF_save_fm DFF_W2467(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D019));
DFF_save_fm DFF_W2468(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D029));
DFF_save_fm DFF_W2469(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D109));
DFF_save_fm DFF_W2470(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D119));
DFF_save_fm DFF_W2471(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D129));
DFF_save_fm DFF_W2472(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D209));
DFF_save_fm DFF_W2473(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D219));
DFF_save_fm DFF_W2474(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D229));
DFF_save_fm DFF_W2475(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D00A));
DFF_save_fm DFF_W2476(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D01A));
DFF_save_fm DFF_W2477(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D02A));
DFF_save_fm DFF_W2478(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D10A));
DFF_save_fm DFF_W2479(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D11A));
DFF_save_fm DFF_W2480(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D12A));
DFF_save_fm DFF_W2481(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D20A));
DFF_save_fm DFF_W2482(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D21A));
DFF_save_fm DFF_W2483(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D22A));
DFF_save_fm DFF_W2484(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D00B));
DFF_save_fm DFF_W2485(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D01B));
DFF_save_fm DFF_W2486(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D02B));
DFF_save_fm DFF_W2487(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D10B));
DFF_save_fm DFF_W2488(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D11B));
DFF_save_fm DFF_W2489(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D12B));
DFF_save_fm DFF_W2490(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D20B));
DFF_save_fm DFF_W2491(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D21B));
DFF_save_fm DFF_W2492(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D22B));
DFF_save_fm DFF_W2493(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D00C));
DFF_save_fm DFF_W2494(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D01C));
DFF_save_fm DFF_W2495(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D02C));
DFF_save_fm DFF_W2496(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D10C));
DFF_save_fm DFF_W2497(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D11C));
DFF_save_fm DFF_W2498(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D12C));
DFF_save_fm DFF_W2499(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D20C));
DFF_save_fm DFF_W2500(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D21C));
DFF_save_fm DFF_W2501(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D22C));
DFF_save_fm DFF_W2502(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D00D));
DFF_save_fm DFF_W2503(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D01D));
DFF_save_fm DFF_W2504(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D02D));
DFF_save_fm DFF_W2505(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D10D));
DFF_save_fm DFF_W2506(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D11D));
DFF_save_fm DFF_W2507(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D12D));
DFF_save_fm DFF_W2508(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D20D));
DFF_save_fm DFF_W2509(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D21D));
DFF_save_fm DFF_W2510(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D22D));
DFF_save_fm DFF_W2511(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D00E));
DFF_save_fm DFF_W2512(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D01E));
DFF_save_fm DFF_W2513(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D02E));
DFF_save_fm DFF_W2514(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D10E));
DFF_save_fm DFF_W2515(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D11E));
DFF_save_fm DFF_W2516(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D12E));
DFF_save_fm DFF_W2517(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D20E));
DFF_save_fm DFF_W2518(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D21E));
DFF_save_fm DFF_W2519(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D22E));
DFF_save_fm DFF_W2520(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D00F));
DFF_save_fm DFF_W2521(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D01F));
DFF_save_fm DFF_W2522(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D02F));
DFF_save_fm DFF_W2523(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D10F));
DFF_save_fm DFF_W2524(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D11F));
DFF_save_fm DFF_W2525(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D12F));
DFF_save_fm DFF_W2526(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D20F));
DFF_save_fm DFF_W2527(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2D21F));
DFF_save_fm DFF_W2528(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2D22F));
DFF_save_fm DFF_W2529(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E000));
DFF_save_fm DFF_W2530(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E010));
DFF_save_fm DFF_W2531(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E020));
DFF_save_fm DFF_W2532(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E100));
DFF_save_fm DFF_W2533(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E110));
DFF_save_fm DFF_W2534(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E120));
DFF_save_fm DFF_W2535(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E200));
DFF_save_fm DFF_W2536(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E210));
DFF_save_fm DFF_W2537(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E220));
DFF_save_fm DFF_W2538(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E001));
DFF_save_fm DFF_W2539(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E011));
DFF_save_fm DFF_W2540(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E021));
DFF_save_fm DFF_W2541(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E101));
DFF_save_fm DFF_W2542(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E111));
DFF_save_fm DFF_W2543(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E121));
DFF_save_fm DFF_W2544(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E201));
DFF_save_fm DFF_W2545(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E211));
DFF_save_fm DFF_W2546(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E221));
DFF_save_fm DFF_W2547(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E002));
DFF_save_fm DFF_W2548(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E012));
DFF_save_fm DFF_W2549(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E022));
DFF_save_fm DFF_W2550(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E102));
DFF_save_fm DFF_W2551(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E112));
DFF_save_fm DFF_W2552(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E122));
DFF_save_fm DFF_W2553(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E202));
DFF_save_fm DFF_W2554(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E212));
DFF_save_fm DFF_W2555(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E222));
DFF_save_fm DFF_W2556(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E003));
DFF_save_fm DFF_W2557(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E013));
DFF_save_fm DFF_W2558(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E023));
DFF_save_fm DFF_W2559(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E103));
DFF_save_fm DFF_W2560(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E113));
DFF_save_fm DFF_W2561(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E123));
DFF_save_fm DFF_W2562(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E203));
DFF_save_fm DFF_W2563(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E213));
DFF_save_fm DFF_W2564(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E223));
DFF_save_fm DFF_W2565(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E004));
DFF_save_fm DFF_W2566(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E014));
DFF_save_fm DFF_W2567(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E024));
DFF_save_fm DFF_W2568(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E104));
DFF_save_fm DFF_W2569(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E114));
DFF_save_fm DFF_W2570(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E124));
DFF_save_fm DFF_W2571(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E204));
DFF_save_fm DFF_W2572(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E214));
DFF_save_fm DFF_W2573(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E224));
DFF_save_fm DFF_W2574(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E005));
DFF_save_fm DFF_W2575(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E015));
DFF_save_fm DFF_W2576(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E025));
DFF_save_fm DFF_W2577(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E105));
DFF_save_fm DFF_W2578(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E115));
DFF_save_fm DFF_W2579(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E125));
DFF_save_fm DFF_W2580(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E205));
DFF_save_fm DFF_W2581(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E215));
DFF_save_fm DFF_W2582(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E225));
DFF_save_fm DFF_W2583(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E006));
DFF_save_fm DFF_W2584(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E016));
DFF_save_fm DFF_W2585(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E026));
DFF_save_fm DFF_W2586(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E106));
DFF_save_fm DFF_W2587(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E116));
DFF_save_fm DFF_W2588(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E126));
DFF_save_fm DFF_W2589(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E206));
DFF_save_fm DFF_W2590(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E216));
DFF_save_fm DFF_W2591(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E226));
DFF_save_fm DFF_W2592(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E007));
DFF_save_fm DFF_W2593(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E017));
DFF_save_fm DFF_W2594(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E027));
DFF_save_fm DFF_W2595(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E107));
DFF_save_fm DFF_W2596(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E117));
DFF_save_fm DFF_W2597(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E127));
DFF_save_fm DFF_W2598(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E207));
DFF_save_fm DFF_W2599(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E217));
DFF_save_fm DFF_W2600(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E227));
DFF_save_fm DFF_W2601(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E008));
DFF_save_fm DFF_W2602(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E018));
DFF_save_fm DFF_W2603(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E028));
DFF_save_fm DFF_W2604(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E108));
DFF_save_fm DFF_W2605(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E118));
DFF_save_fm DFF_W2606(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E128));
DFF_save_fm DFF_W2607(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E208));
DFF_save_fm DFF_W2608(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E218));
DFF_save_fm DFF_W2609(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E228));
DFF_save_fm DFF_W2610(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E009));
DFF_save_fm DFF_W2611(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E019));
DFF_save_fm DFF_W2612(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E029));
DFF_save_fm DFF_W2613(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E109));
DFF_save_fm DFF_W2614(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E119));
DFF_save_fm DFF_W2615(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E129));
DFF_save_fm DFF_W2616(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E209));
DFF_save_fm DFF_W2617(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E219));
DFF_save_fm DFF_W2618(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E229));
DFF_save_fm DFF_W2619(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E00A));
DFF_save_fm DFF_W2620(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E01A));
DFF_save_fm DFF_W2621(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E02A));
DFF_save_fm DFF_W2622(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E10A));
DFF_save_fm DFF_W2623(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E11A));
DFF_save_fm DFF_W2624(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E12A));
DFF_save_fm DFF_W2625(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E20A));
DFF_save_fm DFF_W2626(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E21A));
DFF_save_fm DFF_W2627(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E22A));
DFF_save_fm DFF_W2628(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E00B));
DFF_save_fm DFF_W2629(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E01B));
DFF_save_fm DFF_W2630(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E02B));
DFF_save_fm DFF_W2631(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E10B));
DFF_save_fm DFF_W2632(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E11B));
DFF_save_fm DFF_W2633(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E12B));
DFF_save_fm DFF_W2634(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E20B));
DFF_save_fm DFF_W2635(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E21B));
DFF_save_fm DFF_W2636(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E22B));
DFF_save_fm DFF_W2637(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E00C));
DFF_save_fm DFF_W2638(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E01C));
DFF_save_fm DFF_W2639(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E02C));
DFF_save_fm DFF_W2640(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E10C));
DFF_save_fm DFF_W2641(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E11C));
DFF_save_fm DFF_W2642(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E12C));
DFF_save_fm DFF_W2643(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E20C));
DFF_save_fm DFF_W2644(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E21C));
DFF_save_fm DFF_W2645(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E22C));
DFF_save_fm DFF_W2646(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E00D));
DFF_save_fm DFF_W2647(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E01D));
DFF_save_fm DFF_W2648(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E02D));
DFF_save_fm DFF_W2649(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E10D));
DFF_save_fm DFF_W2650(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E11D));
DFF_save_fm DFF_W2651(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E12D));
DFF_save_fm DFF_W2652(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E20D));
DFF_save_fm DFF_W2653(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E21D));
DFF_save_fm DFF_W2654(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E22D));
DFF_save_fm DFF_W2655(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E00E));
DFF_save_fm DFF_W2656(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E01E));
DFF_save_fm DFF_W2657(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E02E));
DFF_save_fm DFF_W2658(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E10E));
DFF_save_fm DFF_W2659(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E11E));
DFF_save_fm DFF_W2660(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E12E));
DFF_save_fm DFF_W2661(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E20E));
DFF_save_fm DFF_W2662(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E21E));
DFF_save_fm DFF_W2663(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E22E));
DFF_save_fm DFF_W2664(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E00F));
DFF_save_fm DFF_W2665(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E01F));
DFF_save_fm DFF_W2666(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E02F));
DFF_save_fm DFF_W2667(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E10F));
DFF_save_fm DFF_W2668(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E11F));
DFF_save_fm DFF_W2669(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E12F));
DFF_save_fm DFF_W2670(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E20F));
DFF_save_fm DFF_W2671(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2E21F));
DFF_save_fm DFF_W2672(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2E22F));
DFF_save_fm DFF_W2673(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F000));
DFF_save_fm DFF_W2674(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F010));
DFF_save_fm DFF_W2675(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F020));
DFF_save_fm DFF_W2676(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F100));
DFF_save_fm DFF_W2677(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F110));
DFF_save_fm DFF_W2678(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F120));
DFF_save_fm DFF_W2679(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F200));
DFF_save_fm DFF_W2680(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F210));
DFF_save_fm DFF_W2681(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F220));
DFF_save_fm DFF_W2682(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F001));
DFF_save_fm DFF_W2683(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F011));
DFF_save_fm DFF_W2684(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F021));
DFF_save_fm DFF_W2685(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F101));
DFF_save_fm DFF_W2686(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F111));
DFF_save_fm DFF_W2687(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F121));
DFF_save_fm DFF_W2688(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F201));
DFF_save_fm DFF_W2689(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F211));
DFF_save_fm DFF_W2690(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F221));
DFF_save_fm DFF_W2691(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F002));
DFF_save_fm DFF_W2692(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F012));
DFF_save_fm DFF_W2693(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F022));
DFF_save_fm DFF_W2694(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F102));
DFF_save_fm DFF_W2695(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F112));
DFF_save_fm DFF_W2696(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F122));
DFF_save_fm DFF_W2697(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F202));
DFF_save_fm DFF_W2698(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F212));
DFF_save_fm DFF_W2699(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F222));
DFF_save_fm DFF_W2700(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F003));
DFF_save_fm DFF_W2701(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F013));
DFF_save_fm DFF_W2702(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F023));
DFF_save_fm DFF_W2703(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F103));
DFF_save_fm DFF_W2704(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F113));
DFF_save_fm DFF_W2705(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F123));
DFF_save_fm DFF_W2706(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F203));
DFF_save_fm DFF_W2707(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F213));
DFF_save_fm DFF_W2708(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F223));
DFF_save_fm DFF_W2709(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F004));
DFF_save_fm DFF_W2710(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F014));
DFF_save_fm DFF_W2711(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F024));
DFF_save_fm DFF_W2712(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F104));
DFF_save_fm DFF_W2713(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F114));
DFF_save_fm DFF_W2714(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F124));
DFF_save_fm DFF_W2715(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F204));
DFF_save_fm DFF_W2716(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F214));
DFF_save_fm DFF_W2717(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F224));
DFF_save_fm DFF_W2718(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F005));
DFF_save_fm DFF_W2719(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F015));
DFF_save_fm DFF_W2720(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F025));
DFF_save_fm DFF_W2721(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F105));
DFF_save_fm DFF_W2722(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F115));
DFF_save_fm DFF_W2723(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F125));
DFF_save_fm DFF_W2724(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F205));
DFF_save_fm DFF_W2725(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F215));
DFF_save_fm DFF_W2726(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F225));
DFF_save_fm DFF_W2727(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F006));
DFF_save_fm DFF_W2728(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F016));
DFF_save_fm DFF_W2729(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F026));
DFF_save_fm DFF_W2730(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F106));
DFF_save_fm DFF_W2731(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F116));
DFF_save_fm DFF_W2732(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F126));
DFF_save_fm DFF_W2733(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F206));
DFF_save_fm DFF_W2734(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F216));
DFF_save_fm DFF_W2735(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F226));
DFF_save_fm DFF_W2736(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F007));
DFF_save_fm DFF_W2737(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F017));
DFF_save_fm DFF_W2738(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F027));
DFF_save_fm DFF_W2739(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F107));
DFF_save_fm DFF_W2740(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F117));
DFF_save_fm DFF_W2741(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F127));
DFF_save_fm DFF_W2742(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F207));
DFF_save_fm DFF_W2743(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F217));
DFF_save_fm DFF_W2744(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F227));
DFF_save_fm DFF_W2745(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F008));
DFF_save_fm DFF_W2746(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F018));
DFF_save_fm DFF_W2747(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F028));
DFF_save_fm DFF_W2748(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F108));
DFF_save_fm DFF_W2749(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F118));
DFF_save_fm DFF_W2750(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F128));
DFF_save_fm DFF_W2751(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F208));
DFF_save_fm DFF_W2752(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F218));
DFF_save_fm DFF_W2753(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F228));
DFF_save_fm DFF_W2754(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F009));
DFF_save_fm DFF_W2755(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F019));
DFF_save_fm DFF_W2756(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F029));
DFF_save_fm DFF_W2757(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F109));
DFF_save_fm DFF_W2758(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F119));
DFF_save_fm DFF_W2759(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F129));
DFF_save_fm DFF_W2760(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F209));
DFF_save_fm DFF_W2761(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F219));
DFF_save_fm DFF_W2762(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F229));
DFF_save_fm DFF_W2763(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F00A));
DFF_save_fm DFF_W2764(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F01A));
DFF_save_fm DFF_W2765(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F02A));
DFF_save_fm DFF_W2766(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F10A));
DFF_save_fm DFF_W2767(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F11A));
DFF_save_fm DFF_W2768(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F12A));
DFF_save_fm DFF_W2769(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F20A));
DFF_save_fm DFF_W2770(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F21A));
DFF_save_fm DFF_W2771(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F22A));
DFF_save_fm DFF_W2772(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F00B));
DFF_save_fm DFF_W2773(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F01B));
DFF_save_fm DFF_W2774(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F02B));
DFF_save_fm DFF_W2775(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F10B));
DFF_save_fm DFF_W2776(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F11B));
DFF_save_fm DFF_W2777(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F12B));
DFF_save_fm DFF_W2778(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F20B));
DFF_save_fm DFF_W2779(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F21B));
DFF_save_fm DFF_W2780(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F22B));
DFF_save_fm DFF_W2781(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F00C));
DFF_save_fm DFF_W2782(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F01C));
DFF_save_fm DFF_W2783(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F02C));
DFF_save_fm DFF_W2784(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F10C));
DFF_save_fm DFF_W2785(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F11C));
DFF_save_fm DFF_W2786(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F12C));
DFF_save_fm DFF_W2787(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F20C));
DFF_save_fm DFF_W2788(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F21C));
DFF_save_fm DFF_W2789(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F22C));
DFF_save_fm DFF_W2790(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F00D));
DFF_save_fm DFF_W2791(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F01D));
DFF_save_fm DFF_W2792(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F02D));
DFF_save_fm DFF_W2793(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F10D));
DFF_save_fm DFF_W2794(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F11D));
DFF_save_fm DFF_W2795(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F12D));
DFF_save_fm DFF_W2796(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F20D));
DFF_save_fm DFF_W2797(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F21D));
DFF_save_fm DFF_W2798(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F22D));
DFF_save_fm DFF_W2799(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F00E));
DFF_save_fm DFF_W2800(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F01E));
DFF_save_fm DFF_W2801(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F02E));
DFF_save_fm DFF_W2802(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F10E));
DFF_save_fm DFF_W2803(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F11E));
DFF_save_fm DFF_W2804(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F12E));
DFF_save_fm DFF_W2805(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F20E));
DFF_save_fm DFF_W2806(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F21E));
DFF_save_fm DFF_W2807(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F22E));
DFF_save_fm DFF_W2808(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F00F));
DFF_save_fm DFF_W2809(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F01F));
DFF_save_fm DFF_W2810(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F02F));
DFF_save_fm DFF_W2811(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F10F));
DFF_save_fm DFF_W2812(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F11F));
DFF_save_fm DFF_W2813(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F12F));
DFF_save_fm DFF_W2814(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2F20F));
DFF_save_fm DFF_W2815(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F21F));
DFF_save_fm DFF_W2816(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2F22F));
DFF_save_fm DFF_W2817(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G000));
DFF_save_fm DFF_W2818(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G010));
DFF_save_fm DFF_W2819(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G020));
DFF_save_fm DFF_W2820(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G100));
DFF_save_fm DFF_W2821(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G110));
DFF_save_fm DFF_W2822(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G120));
DFF_save_fm DFF_W2823(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G200));
DFF_save_fm DFF_W2824(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G210));
DFF_save_fm DFF_W2825(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G220));
DFF_save_fm DFF_W2826(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G001));
DFF_save_fm DFF_W2827(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G011));
DFF_save_fm DFF_W2828(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G021));
DFF_save_fm DFF_W2829(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G101));
DFF_save_fm DFF_W2830(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G111));
DFF_save_fm DFF_W2831(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G121));
DFF_save_fm DFF_W2832(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G201));
DFF_save_fm DFF_W2833(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G211));
DFF_save_fm DFF_W2834(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G221));
DFF_save_fm DFF_W2835(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G002));
DFF_save_fm DFF_W2836(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G012));
DFF_save_fm DFF_W2837(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G022));
DFF_save_fm DFF_W2838(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G102));
DFF_save_fm DFF_W2839(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G112));
DFF_save_fm DFF_W2840(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G122));
DFF_save_fm DFF_W2841(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G202));
DFF_save_fm DFF_W2842(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G212));
DFF_save_fm DFF_W2843(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G222));
DFF_save_fm DFF_W2844(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G003));
DFF_save_fm DFF_W2845(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G013));
DFF_save_fm DFF_W2846(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G023));
DFF_save_fm DFF_W2847(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G103));
DFF_save_fm DFF_W2848(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G113));
DFF_save_fm DFF_W2849(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G123));
DFF_save_fm DFF_W2850(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G203));
DFF_save_fm DFF_W2851(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G213));
DFF_save_fm DFF_W2852(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G223));
DFF_save_fm DFF_W2853(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G004));
DFF_save_fm DFF_W2854(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G014));
DFF_save_fm DFF_W2855(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G024));
DFF_save_fm DFF_W2856(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G104));
DFF_save_fm DFF_W2857(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G114));
DFF_save_fm DFF_W2858(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G124));
DFF_save_fm DFF_W2859(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G204));
DFF_save_fm DFF_W2860(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G214));
DFF_save_fm DFF_W2861(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G224));
DFF_save_fm DFF_W2862(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G005));
DFF_save_fm DFF_W2863(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G015));
DFF_save_fm DFF_W2864(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G025));
DFF_save_fm DFF_W2865(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G105));
DFF_save_fm DFF_W2866(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G115));
DFF_save_fm DFF_W2867(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G125));
DFF_save_fm DFF_W2868(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G205));
DFF_save_fm DFF_W2869(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G215));
DFF_save_fm DFF_W2870(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G225));
DFF_save_fm DFF_W2871(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G006));
DFF_save_fm DFF_W2872(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G016));
DFF_save_fm DFF_W2873(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G026));
DFF_save_fm DFF_W2874(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G106));
DFF_save_fm DFF_W2875(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G116));
DFF_save_fm DFF_W2876(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G126));
DFF_save_fm DFF_W2877(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G206));
DFF_save_fm DFF_W2878(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G216));
DFF_save_fm DFF_W2879(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G226));
DFF_save_fm DFF_W2880(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G007));
DFF_save_fm DFF_W2881(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G017));
DFF_save_fm DFF_W2882(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G027));
DFF_save_fm DFF_W2883(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G107));
DFF_save_fm DFF_W2884(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G117));
DFF_save_fm DFF_W2885(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G127));
DFF_save_fm DFF_W2886(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G207));
DFF_save_fm DFF_W2887(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G217));
DFF_save_fm DFF_W2888(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G227));
DFF_save_fm DFF_W2889(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G008));
DFF_save_fm DFF_W2890(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G018));
DFF_save_fm DFF_W2891(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G028));
DFF_save_fm DFF_W2892(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G108));
DFF_save_fm DFF_W2893(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G118));
DFF_save_fm DFF_W2894(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G128));
DFF_save_fm DFF_W2895(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G208));
DFF_save_fm DFF_W2896(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G218));
DFF_save_fm DFF_W2897(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G228));
DFF_save_fm DFF_W2898(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G009));
DFF_save_fm DFF_W2899(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G019));
DFF_save_fm DFF_W2900(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G029));
DFF_save_fm DFF_W2901(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G109));
DFF_save_fm DFF_W2902(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G119));
DFF_save_fm DFF_W2903(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G129));
DFF_save_fm DFF_W2904(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G209));
DFF_save_fm DFF_W2905(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G219));
DFF_save_fm DFF_W2906(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G229));
DFF_save_fm DFF_W2907(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G00A));
DFF_save_fm DFF_W2908(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G01A));
DFF_save_fm DFF_W2909(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G02A));
DFF_save_fm DFF_W2910(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G10A));
DFF_save_fm DFF_W2911(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G11A));
DFF_save_fm DFF_W2912(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G12A));
DFF_save_fm DFF_W2913(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G20A));
DFF_save_fm DFF_W2914(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G21A));
DFF_save_fm DFF_W2915(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G22A));
DFF_save_fm DFF_W2916(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G00B));
DFF_save_fm DFF_W2917(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G01B));
DFF_save_fm DFF_W2918(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G02B));
DFF_save_fm DFF_W2919(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G10B));
DFF_save_fm DFF_W2920(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G11B));
DFF_save_fm DFF_W2921(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G12B));
DFF_save_fm DFF_W2922(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G20B));
DFF_save_fm DFF_W2923(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G21B));
DFF_save_fm DFF_W2924(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G22B));
DFF_save_fm DFF_W2925(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G00C));
DFF_save_fm DFF_W2926(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G01C));
DFF_save_fm DFF_W2927(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G02C));
DFF_save_fm DFF_W2928(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G10C));
DFF_save_fm DFF_W2929(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G11C));
DFF_save_fm DFF_W2930(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G12C));
DFF_save_fm DFF_W2931(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G20C));
DFF_save_fm DFF_W2932(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G21C));
DFF_save_fm DFF_W2933(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G22C));
DFF_save_fm DFF_W2934(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G00D));
DFF_save_fm DFF_W2935(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G01D));
DFF_save_fm DFF_W2936(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G02D));
DFF_save_fm DFF_W2937(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G10D));
DFF_save_fm DFF_W2938(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G11D));
DFF_save_fm DFF_W2939(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G12D));
DFF_save_fm DFF_W2940(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G20D));
DFF_save_fm DFF_W2941(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G21D));
DFF_save_fm DFF_W2942(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G22D));
DFF_save_fm DFF_W2943(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G00E));
DFF_save_fm DFF_W2944(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G01E));
DFF_save_fm DFF_W2945(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G02E));
DFF_save_fm DFF_W2946(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G10E));
DFF_save_fm DFF_W2947(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G11E));
DFF_save_fm DFF_W2948(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G12E));
DFF_save_fm DFF_W2949(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G20E));
DFF_save_fm DFF_W2950(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G21E));
DFF_save_fm DFF_W2951(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G22E));
DFF_save_fm DFF_W2952(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G00F));
DFF_save_fm DFF_W2953(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G01F));
DFF_save_fm DFF_W2954(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G02F));
DFF_save_fm DFF_W2955(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G10F));
DFF_save_fm DFF_W2956(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G11F));
DFF_save_fm DFF_W2957(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G12F));
DFF_save_fm DFF_W2958(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2G20F));
DFF_save_fm DFF_W2959(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G21F));
DFF_save_fm DFF_W2960(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2G22F));
DFF_save_fm DFF_W2961(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H000));
DFF_save_fm DFF_W2962(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H010));
DFF_save_fm DFF_W2963(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H020));
DFF_save_fm DFF_W2964(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H100));
DFF_save_fm DFF_W2965(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H110));
DFF_save_fm DFF_W2966(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H120));
DFF_save_fm DFF_W2967(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H200));
DFF_save_fm DFF_W2968(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H210));
DFF_save_fm DFF_W2969(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H220));
DFF_save_fm DFF_W2970(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H001));
DFF_save_fm DFF_W2971(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H011));
DFF_save_fm DFF_W2972(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H021));
DFF_save_fm DFF_W2973(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H101));
DFF_save_fm DFF_W2974(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H111));
DFF_save_fm DFF_W2975(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H121));
DFF_save_fm DFF_W2976(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H201));
DFF_save_fm DFF_W2977(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H211));
DFF_save_fm DFF_W2978(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H221));
DFF_save_fm DFF_W2979(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H002));
DFF_save_fm DFF_W2980(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H012));
DFF_save_fm DFF_W2981(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H022));
DFF_save_fm DFF_W2982(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H102));
DFF_save_fm DFF_W2983(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H112));
DFF_save_fm DFF_W2984(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H122));
DFF_save_fm DFF_W2985(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H202));
DFF_save_fm DFF_W2986(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H212));
DFF_save_fm DFF_W2987(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H222));
DFF_save_fm DFF_W2988(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H003));
DFF_save_fm DFF_W2989(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H013));
DFF_save_fm DFF_W2990(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H023));
DFF_save_fm DFF_W2991(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H103));
DFF_save_fm DFF_W2992(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H113));
DFF_save_fm DFF_W2993(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H123));
DFF_save_fm DFF_W2994(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H203));
DFF_save_fm DFF_W2995(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H213));
DFF_save_fm DFF_W2996(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H223));
DFF_save_fm DFF_W2997(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H004));
DFF_save_fm DFF_W2998(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H014));
DFF_save_fm DFF_W2999(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H024));
DFF_save_fm DFF_W3000(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H104));
DFF_save_fm DFF_W3001(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H114));
DFF_save_fm DFF_W3002(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H124));
DFF_save_fm DFF_W3003(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H204));
DFF_save_fm DFF_W3004(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H214));
DFF_save_fm DFF_W3005(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H224));
DFF_save_fm DFF_W3006(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H005));
DFF_save_fm DFF_W3007(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H015));
DFF_save_fm DFF_W3008(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H025));
DFF_save_fm DFF_W3009(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H105));
DFF_save_fm DFF_W3010(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H115));
DFF_save_fm DFF_W3011(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H125));
DFF_save_fm DFF_W3012(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H205));
DFF_save_fm DFF_W3013(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H215));
DFF_save_fm DFF_W3014(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H225));
DFF_save_fm DFF_W3015(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H006));
DFF_save_fm DFF_W3016(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H016));
DFF_save_fm DFF_W3017(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H026));
DFF_save_fm DFF_W3018(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H106));
DFF_save_fm DFF_W3019(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H116));
DFF_save_fm DFF_W3020(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H126));
DFF_save_fm DFF_W3021(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H206));
DFF_save_fm DFF_W3022(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H216));
DFF_save_fm DFF_W3023(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H226));
DFF_save_fm DFF_W3024(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H007));
DFF_save_fm DFF_W3025(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H017));
DFF_save_fm DFF_W3026(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H027));
DFF_save_fm DFF_W3027(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H107));
DFF_save_fm DFF_W3028(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H117));
DFF_save_fm DFF_W3029(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H127));
DFF_save_fm DFF_W3030(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H207));
DFF_save_fm DFF_W3031(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H217));
DFF_save_fm DFF_W3032(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H227));
DFF_save_fm DFF_W3033(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H008));
DFF_save_fm DFF_W3034(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H018));
DFF_save_fm DFF_W3035(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H028));
DFF_save_fm DFF_W3036(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H108));
DFF_save_fm DFF_W3037(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H118));
DFF_save_fm DFF_W3038(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H128));
DFF_save_fm DFF_W3039(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H208));
DFF_save_fm DFF_W3040(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H218));
DFF_save_fm DFF_W3041(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H228));
DFF_save_fm DFF_W3042(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H009));
DFF_save_fm DFF_W3043(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H019));
DFF_save_fm DFF_W3044(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H029));
DFF_save_fm DFF_W3045(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H109));
DFF_save_fm DFF_W3046(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H119));
DFF_save_fm DFF_W3047(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H129));
DFF_save_fm DFF_W3048(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H209));
DFF_save_fm DFF_W3049(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H219));
DFF_save_fm DFF_W3050(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H229));
DFF_save_fm DFF_W3051(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H00A));
DFF_save_fm DFF_W3052(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H01A));
DFF_save_fm DFF_W3053(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H02A));
DFF_save_fm DFF_W3054(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H10A));
DFF_save_fm DFF_W3055(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H11A));
DFF_save_fm DFF_W3056(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H12A));
DFF_save_fm DFF_W3057(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H20A));
DFF_save_fm DFF_W3058(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H21A));
DFF_save_fm DFF_W3059(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H22A));
DFF_save_fm DFF_W3060(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H00B));
DFF_save_fm DFF_W3061(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H01B));
DFF_save_fm DFF_W3062(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H02B));
DFF_save_fm DFF_W3063(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H10B));
DFF_save_fm DFF_W3064(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H11B));
DFF_save_fm DFF_W3065(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H12B));
DFF_save_fm DFF_W3066(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H20B));
DFF_save_fm DFF_W3067(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H21B));
DFF_save_fm DFF_W3068(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H22B));
DFF_save_fm DFF_W3069(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H00C));
DFF_save_fm DFF_W3070(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H01C));
DFF_save_fm DFF_W3071(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H02C));
DFF_save_fm DFF_W3072(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H10C));
DFF_save_fm DFF_W3073(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H11C));
DFF_save_fm DFF_W3074(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H12C));
DFF_save_fm DFF_W3075(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H20C));
DFF_save_fm DFF_W3076(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H21C));
DFF_save_fm DFF_W3077(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H22C));
DFF_save_fm DFF_W3078(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H00D));
DFF_save_fm DFF_W3079(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H01D));
DFF_save_fm DFF_W3080(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H02D));
DFF_save_fm DFF_W3081(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H10D));
DFF_save_fm DFF_W3082(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H11D));
DFF_save_fm DFF_W3083(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H12D));
DFF_save_fm DFF_W3084(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H20D));
DFF_save_fm DFF_W3085(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H21D));
DFF_save_fm DFF_W3086(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H22D));
DFF_save_fm DFF_W3087(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H00E));
DFF_save_fm DFF_W3088(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H01E));
DFF_save_fm DFF_W3089(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H02E));
DFF_save_fm DFF_W3090(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H10E));
DFF_save_fm DFF_W3091(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H11E));
DFF_save_fm DFF_W3092(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H12E));
DFF_save_fm DFF_W3093(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H20E));
DFF_save_fm DFF_W3094(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H21E));
DFF_save_fm DFF_W3095(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H22E));
DFF_save_fm DFF_W3096(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H00F));
DFF_save_fm DFF_W3097(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H01F));
DFF_save_fm DFF_W3098(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H02F));
DFF_save_fm DFF_W3099(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H10F));
DFF_save_fm DFF_W3100(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H11F));
DFF_save_fm DFF_W3101(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H12F));
DFF_save_fm DFF_W3102(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H20F));
DFF_save_fm DFF_W3103(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2H21F));
DFF_save_fm DFF_W3104(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2H22F));
DFF_save_fm DFF_W3105(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I000));
DFF_save_fm DFF_W3106(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I010));
DFF_save_fm DFF_W3107(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I020));
DFF_save_fm DFF_W3108(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I100));
DFF_save_fm DFF_W3109(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I110));
DFF_save_fm DFF_W3110(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I120));
DFF_save_fm DFF_W3111(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I200));
DFF_save_fm DFF_W3112(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I210));
DFF_save_fm DFF_W3113(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I220));
DFF_save_fm DFF_W3114(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I001));
DFF_save_fm DFF_W3115(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I011));
DFF_save_fm DFF_W3116(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I021));
DFF_save_fm DFF_W3117(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I101));
DFF_save_fm DFF_W3118(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I111));
DFF_save_fm DFF_W3119(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I121));
DFF_save_fm DFF_W3120(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I201));
DFF_save_fm DFF_W3121(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I211));
DFF_save_fm DFF_W3122(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I221));
DFF_save_fm DFF_W3123(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I002));
DFF_save_fm DFF_W3124(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I012));
DFF_save_fm DFF_W3125(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I022));
DFF_save_fm DFF_W3126(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I102));
DFF_save_fm DFF_W3127(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I112));
DFF_save_fm DFF_W3128(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I122));
DFF_save_fm DFF_W3129(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I202));
DFF_save_fm DFF_W3130(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I212));
DFF_save_fm DFF_W3131(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I222));
DFF_save_fm DFF_W3132(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I003));
DFF_save_fm DFF_W3133(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I013));
DFF_save_fm DFF_W3134(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I023));
DFF_save_fm DFF_W3135(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I103));
DFF_save_fm DFF_W3136(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I113));
DFF_save_fm DFF_W3137(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I123));
DFF_save_fm DFF_W3138(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I203));
DFF_save_fm DFF_W3139(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I213));
DFF_save_fm DFF_W3140(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I223));
DFF_save_fm DFF_W3141(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I004));
DFF_save_fm DFF_W3142(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I014));
DFF_save_fm DFF_W3143(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I024));
DFF_save_fm DFF_W3144(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I104));
DFF_save_fm DFF_W3145(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I114));
DFF_save_fm DFF_W3146(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I124));
DFF_save_fm DFF_W3147(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I204));
DFF_save_fm DFF_W3148(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I214));
DFF_save_fm DFF_W3149(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I224));
DFF_save_fm DFF_W3150(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I005));
DFF_save_fm DFF_W3151(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I015));
DFF_save_fm DFF_W3152(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I025));
DFF_save_fm DFF_W3153(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I105));
DFF_save_fm DFF_W3154(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I115));
DFF_save_fm DFF_W3155(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I125));
DFF_save_fm DFF_W3156(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I205));
DFF_save_fm DFF_W3157(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I215));
DFF_save_fm DFF_W3158(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I225));
DFF_save_fm DFF_W3159(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I006));
DFF_save_fm DFF_W3160(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I016));
DFF_save_fm DFF_W3161(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I026));
DFF_save_fm DFF_W3162(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I106));
DFF_save_fm DFF_W3163(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I116));
DFF_save_fm DFF_W3164(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I126));
DFF_save_fm DFF_W3165(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I206));
DFF_save_fm DFF_W3166(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I216));
DFF_save_fm DFF_W3167(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I226));
DFF_save_fm DFF_W3168(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I007));
DFF_save_fm DFF_W3169(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I017));
DFF_save_fm DFF_W3170(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I027));
DFF_save_fm DFF_W3171(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I107));
DFF_save_fm DFF_W3172(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I117));
DFF_save_fm DFF_W3173(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I127));
DFF_save_fm DFF_W3174(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I207));
DFF_save_fm DFF_W3175(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I217));
DFF_save_fm DFF_W3176(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I227));
DFF_save_fm DFF_W3177(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I008));
DFF_save_fm DFF_W3178(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I018));
DFF_save_fm DFF_W3179(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I028));
DFF_save_fm DFF_W3180(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I108));
DFF_save_fm DFF_W3181(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I118));
DFF_save_fm DFF_W3182(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I128));
DFF_save_fm DFF_W3183(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I208));
DFF_save_fm DFF_W3184(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I218));
DFF_save_fm DFF_W3185(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I228));
DFF_save_fm DFF_W3186(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I009));
DFF_save_fm DFF_W3187(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I019));
DFF_save_fm DFF_W3188(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I029));
DFF_save_fm DFF_W3189(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I109));
DFF_save_fm DFF_W3190(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I119));
DFF_save_fm DFF_W3191(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I129));
DFF_save_fm DFF_W3192(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I209));
DFF_save_fm DFF_W3193(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I219));
DFF_save_fm DFF_W3194(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I229));
DFF_save_fm DFF_W3195(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I00A));
DFF_save_fm DFF_W3196(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I01A));
DFF_save_fm DFF_W3197(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I02A));
DFF_save_fm DFF_W3198(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I10A));
DFF_save_fm DFF_W3199(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I11A));
DFF_save_fm DFF_W3200(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I12A));
DFF_save_fm DFF_W3201(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I20A));
DFF_save_fm DFF_W3202(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I21A));
DFF_save_fm DFF_W3203(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I22A));
DFF_save_fm DFF_W3204(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I00B));
DFF_save_fm DFF_W3205(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I01B));
DFF_save_fm DFF_W3206(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I02B));
DFF_save_fm DFF_W3207(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I10B));
DFF_save_fm DFF_W3208(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I11B));
DFF_save_fm DFF_W3209(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I12B));
DFF_save_fm DFF_W3210(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I20B));
DFF_save_fm DFF_W3211(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I21B));
DFF_save_fm DFF_W3212(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I22B));
DFF_save_fm DFF_W3213(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I00C));
DFF_save_fm DFF_W3214(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I01C));
DFF_save_fm DFF_W3215(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I02C));
DFF_save_fm DFF_W3216(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I10C));
DFF_save_fm DFF_W3217(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I11C));
DFF_save_fm DFF_W3218(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I12C));
DFF_save_fm DFF_W3219(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I20C));
DFF_save_fm DFF_W3220(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I21C));
DFF_save_fm DFF_W3221(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I22C));
DFF_save_fm DFF_W3222(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I00D));
DFF_save_fm DFF_W3223(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I01D));
DFF_save_fm DFF_W3224(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I02D));
DFF_save_fm DFF_W3225(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I10D));
DFF_save_fm DFF_W3226(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I11D));
DFF_save_fm DFF_W3227(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I12D));
DFF_save_fm DFF_W3228(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I20D));
DFF_save_fm DFF_W3229(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I21D));
DFF_save_fm DFF_W3230(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I22D));
DFF_save_fm DFF_W3231(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I00E));
DFF_save_fm DFF_W3232(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I01E));
DFF_save_fm DFF_W3233(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I02E));
DFF_save_fm DFF_W3234(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I10E));
DFF_save_fm DFF_W3235(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I11E));
DFF_save_fm DFF_W3236(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I12E));
DFF_save_fm DFF_W3237(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I20E));
DFF_save_fm DFF_W3238(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I21E));
DFF_save_fm DFF_W3239(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I22E));
DFF_save_fm DFF_W3240(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I00F));
DFF_save_fm DFF_W3241(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I01F));
DFF_save_fm DFF_W3242(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I02F));
DFF_save_fm DFF_W3243(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I10F));
DFF_save_fm DFF_W3244(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I11F));
DFF_save_fm DFF_W3245(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I12F));
DFF_save_fm DFF_W3246(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I20F));
DFF_save_fm DFF_W3247(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2I21F));
DFF_save_fm DFF_W3248(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2I22F));
DFF_save_fm DFF_W3249(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J000));
DFF_save_fm DFF_W3250(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J010));
DFF_save_fm DFF_W3251(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J020));
DFF_save_fm DFF_W3252(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J100));
DFF_save_fm DFF_W3253(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J110));
DFF_save_fm DFF_W3254(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J120));
DFF_save_fm DFF_W3255(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J200));
DFF_save_fm DFF_W3256(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J210));
DFF_save_fm DFF_W3257(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J220));
DFF_save_fm DFF_W3258(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J001));
DFF_save_fm DFF_W3259(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J011));
DFF_save_fm DFF_W3260(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J021));
DFF_save_fm DFF_W3261(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J101));
DFF_save_fm DFF_W3262(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J111));
DFF_save_fm DFF_W3263(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J121));
DFF_save_fm DFF_W3264(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J201));
DFF_save_fm DFF_W3265(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J211));
DFF_save_fm DFF_W3266(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J221));
DFF_save_fm DFF_W3267(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J002));
DFF_save_fm DFF_W3268(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J012));
DFF_save_fm DFF_W3269(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J022));
DFF_save_fm DFF_W3270(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J102));
DFF_save_fm DFF_W3271(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J112));
DFF_save_fm DFF_W3272(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J122));
DFF_save_fm DFF_W3273(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J202));
DFF_save_fm DFF_W3274(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J212));
DFF_save_fm DFF_W3275(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J222));
DFF_save_fm DFF_W3276(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J003));
DFF_save_fm DFF_W3277(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J013));
DFF_save_fm DFF_W3278(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J023));
DFF_save_fm DFF_W3279(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J103));
DFF_save_fm DFF_W3280(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J113));
DFF_save_fm DFF_W3281(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J123));
DFF_save_fm DFF_W3282(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J203));
DFF_save_fm DFF_W3283(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J213));
DFF_save_fm DFF_W3284(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J223));
DFF_save_fm DFF_W3285(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J004));
DFF_save_fm DFF_W3286(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J014));
DFF_save_fm DFF_W3287(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J024));
DFF_save_fm DFF_W3288(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J104));
DFF_save_fm DFF_W3289(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J114));
DFF_save_fm DFF_W3290(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J124));
DFF_save_fm DFF_W3291(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J204));
DFF_save_fm DFF_W3292(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J214));
DFF_save_fm DFF_W3293(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J224));
DFF_save_fm DFF_W3294(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J005));
DFF_save_fm DFF_W3295(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J015));
DFF_save_fm DFF_W3296(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J025));
DFF_save_fm DFF_W3297(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J105));
DFF_save_fm DFF_W3298(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J115));
DFF_save_fm DFF_W3299(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J125));
DFF_save_fm DFF_W3300(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J205));
DFF_save_fm DFF_W3301(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J215));
DFF_save_fm DFF_W3302(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J225));
DFF_save_fm DFF_W3303(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J006));
DFF_save_fm DFF_W3304(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J016));
DFF_save_fm DFF_W3305(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J026));
DFF_save_fm DFF_W3306(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J106));
DFF_save_fm DFF_W3307(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J116));
DFF_save_fm DFF_W3308(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J126));
DFF_save_fm DFF_W3309(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J206));
DFF_save_fm DFF_W3310(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J216));
DFF_save_fm DFF_W3311(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J226));
DFF_save_fm DFF_W3312(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J007));
DFF_save_fm DFF_W3313(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J017));
DFF_save_fm DFF_W3314(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J027));
DFF_save_fm DFF_W3315(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J107));
DFF_save_fm DFF_W3316(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J117));
DFF_save_fm DFF_W3317(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J127));
DFF_save_fm DFF_W3318(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J207));
DFF_save_fm DFF_W3319(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J217));
DFF_save_fm DFF_W3320(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J227));
DFF_save_fm DFF_W3321(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J008));
DFF_save_fm DFF_W3322(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J018));
DFF_save_fm DFF_W3323(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J028));
DFF_save_fm DFF_W3324(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J108));
DFF_save_fm DFF_W3325(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J118));
DFF_save_fm DFF_W3326(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J128));
DFF_save_fm DFF_W3327(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J208));
DFF_save_fm DFF_W3328(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J218));
DFF_save_fm DFF_W3329(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J228));
DFF_save_fm DFF_W3330(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J009));
DFF_save_fm DFF_W3331(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J019));
DFF_save_fm DFF_W3332(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J029));
DFF_save_fm DFF_W3333(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J109));
DFF_save_fm DFF_W3334(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J119));
DFF_save_fm DFF_W3335(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J129));
DFF_save_fm DFF_W3336(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J209));
DFF_save_fm DFF_W3337(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J219));
DFF_save_fm DFF_W3338(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J229));
DFF_save_fm DFF_W3339(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J00A));
DFF_save_fm DFF_W3340(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J01A));
DFF_save_fm DFF_W3341(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J02A));
DFF_save_fm DFF_W3342(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J10A));
DFF_save_fm DFF_W3343(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J11A));
DFF_save_fm DFF_W3344(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J12A));
DFF_save_fm DFF_W3345(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J20A));
DFF_save_fm DFF_W3346(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J21A));
DFF_save_fm DFF_W3347(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J22A));
DFF_save_fm DFF_W3348(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J00B));
DFF_save_fm DFF_W3349(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J01B));
DFF_save_fm DFF_W3350(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J02B));
DFF_save_fm DFF_W3351(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J10B));
DFF_save_fm DFF_W3352(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J11B));
DFF_save_fm DFF_W3353(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J12B));
DFF_save_fm DFF_W3354(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J20B));
DFF_save_fm DFF_W3355(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J21B));
DFF_save_fm DFF_W3356(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J22B));
DFF_save_fm DFF_W3357(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J00C));
DFF_save_fm DFF_W3358(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J01C));
DFF_save_fm DFF_W3359(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J02C));
DFF_save_fm DFF_W3360(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J10C));
DFF_save_fm DFF_W3361(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J11C));
DFF_save_fm DFF_W3362(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J12C));
DFF_save_fm DFF_W3363(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J20C));
DFF_save_fm DFF_W3364(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J21C));
DFF_save_fm DFF_W3365(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J22C));
DFF_save_fm DFF_W3366(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J00D));
DFF_save_fm DFF_W3367(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J01D));
DFF_save_fm DFF_W3368(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J02D));
DFF_save_fm DFF_W3369(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J10D));
DFF_save_fm DFF_W3370(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J11D));
DFF_save_fm DFF_W3371(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J12D));
DFF_save_fm DFF_W3372(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J20D));
DFF_save_fm DFF_W3373(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J21D));
DFF_save_fm DFF_W3374(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J22D));
DFF_save_fm DFF_W3375(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J00E));
DFF_save_fm DFF_W3376(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J01E));
DFF_save_fm DFF_W3377(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J02E));
DFF_save_fm DFF_W3378(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J10E));
DFF_save_fm DFF_W3379(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J11E));
DFF_save_fm DFF_W3380(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J12E));
DFF_save_fm DFF_W3381(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J20E));
DFF_save_fm DFF_W3382(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J21E));
DFF_save_fm DFF_W3383(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J22E));
DFF_save_fm DFF_W3384(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J00F));
DFF_save_fm DFF_W3385(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2J01F));
DFF_save_fm DFF_W3386(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J02F));
DFF_save_fm DFF_W3387(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J10F));
DFF_save_fm DFF_W3388(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J11F));
DFF_save_fm DFF_W3389(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J12F));
DFF_save_fm DFF_W3390(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J20F));
DFF_save_fm DFF_W3391(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J21F));
DFF_save_fm DFF_W3392(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2J22F));
DFF_save_fm DFF_W3393(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K000));
DFF_save_fm DFF_W3394(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K010));
DFF_save_fm DFF_W3395(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K020));
DFF_save_fm DFF_W3396(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K100));
DFF_save_fm DFF_W3397(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K110));
DFF_save_fm DFF_W3398(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K120));
DFF_save_fm DFF_W3399(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K200));
DFF_save_fm DFF_W3400(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K210));
DFF_save_fm DFF_W3401(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K220));
DFF_save_fm DFF_W3402(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K001));
DFF_save_fm DFF_W3403(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K011));
DFF_save_fm DFF_W3404(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K021));
DFF_save_fm DFF_W3405(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K101));
DFF_save_fm DFF_W3406(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K111));
DFF_save_fm DFF_W3407(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K121));
DFF_save_fm DFF_W3408(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K201));
DFF_save_fm DFF_W3409(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K211));
DFF_save_fm DFF_W3410(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K221));
DFF_save_fm DFF_W3411(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K002));
DFF_save_fm DFF_W3412(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K012));
DFF_save_fm DFF_W3413(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K022));
DFF_save_fm DFF_W3414(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K102));
DFF_save_fm DFF_W3415(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K112));
DFF_save_fm DFF_W3416(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K122));
DFF_save_fm DFF_W3417(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K202));
DFF_save_fm DFF_W3418(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K212));
DFF_save_fm DFF_W3419(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K222));
DFF_save_fm DFF_W3420(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K003));
DFF_save_fm DFF_W3421(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K013));
DFF_save_fm DFF_W3422(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K023));
DFF_save_fm DFF_W3423(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K103));
DFF_save_fm DFF_W3424(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K113));
DFF_save_fm DFF_W3425(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K123));
DFF_save_fm DFF_W3426(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K203));
DFF_save_fm DFF_W3427(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K213));
DFF_save_fm DFF_W3428(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K223));
DFF_save_fm DFF_W3429(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K004));
DFF_save_fm DFF_W3430(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K014));
DFF_save_fm DFF_W3431(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K024));
DFF_save_fm DFF_W3432(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K104));
DFF_save_fm DFF_W3433(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K114));
DFF_save_fm DFF_W3434(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K124));
DFF_save_fm DFF_W3435(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K204));
DFF_save_fm DFF_W3436(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K214));
DFF_save_fm DFF_W3437(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K224));
DFF_save_fm DFF_W3438(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K005));
DFF_save_fm DFF_W3439(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K015));
DFF_save_fm DFF_W3440(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K025));
DFF_save_fm DFF_W3441(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K105));
DFF_save_fm DFF_W3442(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K115));
DFF_save_fm DFF_W3443(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K125));
DFF_save_fm DFF_W3444(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K205));
DFF_save_fm DFF_W3445(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K215));
DFF_save_fm DFF_W3446(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K225));
DFF_save_fm DFF_W3447(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K006));
DFF_save_fm DFF_W3448(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K016));
DFF_save_fm DFF_W3449(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K026));
DFF_save_fm DFF_W3450(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K106));
DFF_save_fm DFF_W3451(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K116));
DFF_save_fm DFF_W3452(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K126));
DFF_save_fm DFF_W3453(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K206));
DFF_save_fm DFF_W3454(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K216));
DFF_save_fm DFF_W3455(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K226));
DFF_save_fm DFF_W3456(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K007));
DFF_save_fm DFF_W3457(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K017));
DFF_save_fm DFF_W3458(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K027));
DFF_save_fm DFF_W3459(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K107));
DFF_save_fm DFF_W3460(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K117));
DFF_save_fm DFF_W3461(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K127));
DFF_save_fm DFF_W3462(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K207));
DFF_save_fm DFF_W3463(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K217));
DFF_save_fm DFF_W3464(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K227));
DFF_save_fm DFF_W3465(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K008));
DFF_save_fm DFF_W3466(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K018));
DFF_save_fm DFF_W3467(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K028));
DFF_save_fm DFF_W3468(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K108));
DFF_save_fm DFF_W3469(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K118));
DFF_save_fm DFF_W3470(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K128));
DFF_save_fm DFF_W3471(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K208));
DFF_save_fm DFF_W3472(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K218));
DFF_save_fm DFF_W3473(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K228));
DFF_save_fm DFF_W3474(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K009));
DFF_save_fm DFF_W3475(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K019));
DFF_save_fm DFF_W3476(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K029));
DFF_save_fm DFF_W3477(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K109));
DFF_save_fm DFF_W3478(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K119));
DFF_save_fm DFF_W3479(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K129));
DFF_save_fm DFF_W3480(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K209));
DFF_save_fm DFF_W3481(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K219));
DFF_save_fm DFF_W3482(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K229));
DFF_save_fm DFF_W3483(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K00A));
DFF_save_fm DFF_W3484(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K01A));
DFF_save_fm DFF_W3485(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K02A));
DFF_save_fm DFF_W3486(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K10A));
DFF_save_fm DFF_W3487(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K11A));
DFF_save_fm DFF_W3488(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K12A));
DFF_save_fm DFF_W3489(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K20A));
DFF_save_fm DFF_W3490(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K21A));
DFF_save_fm DFF_W3491(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K22A));
DFF_save_fm DFF_W3492(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K00B));
DFF_save_fm DFF_W3493(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K01B));
DFF_save_fm DFF_W3494(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K02B));
DFF_save_fm DFF_W3495(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K10B));
DFF_save_fm DFF_W3496(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K11B));
DFF_save_fm DFF_W3497(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K12B));
DFF_save_fm DFF_W3498(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K20B));
DFF_save_fm DFF_W3499(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K21B));
DFF_save_fm DFF_W3500(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K22B));
DFF_save_fm DFF_W3501(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K00C));
DFF_save_fm DFF_W3502(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K01C));
DFF_save_fm DFF_W3503(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K02C));
DFF_save_fm DFF_W3504(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K10C));
DFF_save_fm DFF_W3505(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K11C));
DFF_save_fm DFF_W3506(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K12C));
DFF_save_fm DFF_W3507(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K20C));
DFF_save_fm DFF_W3508(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K21C));
DFF_save_fm DFF_W3509(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K22C));
DFF_save_fm DFF_W3510(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K00D));
DFF_save_fm DFF_W3511(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K01D));
DFF_save_fm DFF_W3512(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K02D));
DFF_save_fm DFF_W3513(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K10D));
DFF_save_fm DFF_W3514(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K11D));
DFF_save_fm DFF_W3515(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K12D));
DFF_save_fm DFF_W3516(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K20D));
DFF_save_fm DFF_W3517(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K21D));
DFF_save_fm DFF_W3518(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K22D));
DFF_save_fm DFF_W3519(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K00E));
DFF_save_fm DFF_W3520(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K01E));
DFF_save_fm DFF_W3521(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K02E));
DFF_save_fm DFF_W3522(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K10E));
DFF_save_fm DFF_W3523(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K11E));
DFF_save_fm DFF_W3524(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K12E));
DFF_save_fm DFF_W3525(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K20E));
DFF_save_fm DFF_W3526(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K21E));
DFF_save_fm DFF_W3527(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K22E));
DFF_save_fm DFF_W3528(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K00F));
DFF_save_fm DFF_W3529(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K01F));
DFF_save_fm DFF_W3530(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K02F));
DFF_save_fm DFF_W3531(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K10F));
DFF_save_fm DFF_W3532(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K11F));
DFF_save_fm DFF_W3533(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K12F));
DFF_save_fm DFF_W3534(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K20F));
DFF_save_fm DFF_W3535(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2K21F));
DFF_save_fm DFF_W3536(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2K22F));
DFF_save_fm DFF_W3537(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L000));
DFF_save_fm DFF_W3538(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L010));
DFF_save_fm DFF_W3539(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L020));
DFF_save_fm DFF_W3540(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L100));
DFF_save_fm DFF_W3541(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L110));
DFF_save_fm DFF_W3542(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L120));
DFF_save_fm DFF_W3543(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L200));
DFF_save_fm DFF_W3544(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L210));
DFF_save_fm DFF_W3545(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L220));
DFF_save_fm DFF_W3546(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L001));
DFF_save_fm DFF_W3547(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L011));
DFF_save_fm DFF_W3548(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L021));
DFF_save_fm DFF_W3549(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L101));
DFF_save_fm DFF_W3550(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L111));
DFF_save_fm DFF_W3551(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L121));
DFF_save_fm DFF_W3552(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L201));
DFF_save_fm DFF_W3553(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L211));
DFF_save_fm DFF_W3554(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L221));
DFF_save_fm DFF_W3555(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L002));
DFF_save_fm DFF_W3556(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L012));
DFF_save_fm DFF_W3557(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L022));
DFF_save_fm DFF_W3558(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L102));
DFF_save_fm DFF_W3559(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L112));
DFF_save_fm DFF_W3560(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L122));
DFF_save_fm DFF_W3561(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L202));
DFF_save_fm DFF_W3562(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L212));
DFF_save_fm DFF_W3563(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L222));
DFF_save_fm DFF_W3564(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L003));
DFF_save_fm DFF_W3565(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L013));
DFF_save_fm DFF_W3566(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L023));
DFF_save_fm DFF_W3567(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L103));
DFF_save_fm DFF_W3568(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L113));
DFF_save_fm DFF_W3569(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L123));
DFF_save_fm DFF_W3570(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L203));
DFF_save_fm DFF_W3571(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L213));
DFF_save_fm DFF_W3572(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L223));
DFF_save_fm DFF_W3573(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L004));
DFF_save_fm DFF_W3574(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L014));
DFF_save_fm DFF_W3575(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L024));
DFF_save_fm DFF_W3576(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L104));
DFF_save_fm DFF_W3577(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L114));
DFF_save_fm DFF_W3578(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L124));
DFF_save_fm DFF_W3579(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L204));
DFF_save_fm DFF_W3580(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L214));
DFF_save_fm DFF_W3581(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L224));
DFF_save_fm DFF_W3582(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L005));
DFF_save_fm DFF_W3583(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L015));
DFF_save_fm DFF_W3584(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L025));
DFF_save_fm DFF_W3585(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L105));
DFF_save_fm DFF_W3586(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L115));
DFF_save_fm DFF_W3587(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L125));
DFF_save_fm DFF_W3588(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L205));
DFF_save_fm DFF_W3589(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L215));
DFF_save_fm DFF_W3590(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L225));
DFF_save_fm DFF_W3591(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L006));
DFF_save_fm DFF_W3592(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L016));
DFF_save_fm DFF_W3593(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L026));
DFF_save_fm DFF_W3594(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L106));
DFF_save_fm DFF_W3595(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L116));
DFF_save_fm DFF_W3596(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L126));
DFF_save_fm DFF_W3597(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L206));
DFF_save_fm DFF_W3598(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L216));
DFF_save_fm DFF_W3599(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L226));
DFF_save_fm DFF_W3600(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L007));
DFF_save_fm DFF_W3601(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L017));
DFF_save_fm DFF_W3602(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L027));
DFF_save_fm DFF_W3603(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L107));
DFF_save_fm DFF_W3604(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L117));
DFF_save_fm DFF_W3605(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L127));
DFF_save_fm DFF_W3606(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L207));
DFF_save_fm DFF_W3607(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L217));
DFF_save_fm DFF_W3608(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L227));
DFF_save_fm DFF_W3609(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L008));
DFF_save_fm DFF_W3610(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L018));
DFF_save_fm DFF_W3611(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L028));
DFF_save_fm DFF_W3612(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L108));
DFF_save_fm DFF_W3613(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L118));
DFF_save_fm DFF_W3614(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L128));
DFF_save_fm DFF_W3615(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L208));
DFF_save_fm DFF_W3616(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L218));
DFF_save_fm DFF_W3617(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L228));
DFF_save_fm DFF_W3618(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L009));
DFF_save_fm DFF_W3619(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L019));
DFF_save_fm DFF_W3620(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L029));
DFF_save_fm DFF_W3621(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L109));
DFF_save_fm DFF_W3622(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L119));
DFF_save_fm DFF_W3623(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L129));
DFF_save_fm DFF_W3624(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L209));
DFF_save_fm DFF_W3625(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L219));
DFF_save_fm DFF_W3626(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L229));
DFF_save_fm DFF_W3627(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L00A));
DFF_save_fm DFF_W3628(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L01A));
DFF_save_fm DFF_W3629(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L02A));
DFF_save_fm DFF_W3630(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L10A));
DFF_save_fm DFF_W3631(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L11A));
DFF_save_fm DFF_W3632(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L12A));
DFF_save_fm DFF_W3633(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L20A));
DFF_save_fm DFF_W3634(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L21A));
DFF_save_fm DFF_W3635(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L22A));
DFF_save_fm DFF_W3636(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L00B));
DFF_save_fm DFF_W3637(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L01B));
DFF_save_fm DFF_W3638(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L02B));
DFF_save_fm DFF_W3639(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L10B));
DFF_save_fm DFF_W3640(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L11B));
DFF_save_fm DFF_W3641(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L12B));
DFF_save_fm DFF_W3642(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L20B));
DFF_save_fm DFF_W3643(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L21B));
DFF_save_fm DFF_W3644(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L22B));
DFF_save_fm DFF_W3645(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L00C));
DFF_save_fm DFF_W3646(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L01C));
DFF_save_fm DFF_W3647(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L02C));
DFF_save_fm DFF_W3648(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L10C));
DFF_save_fm DFF_W3649(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L11C));
DFF_save_fm DFF_W3650(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L12C));
DFF_save_fm DFF_W3651(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L20C));
DFF_save_fm DFF_W3652(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L21C));
DFF_save_fm DFF_W3653(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L22C));
DFF_save_fm DFF_W3654(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L00D));
DFF_save_fm DFF_W3655(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L01D));
DFF_save_fm DFF_W3656(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L02D));
DFF_save_fm DFF_W3657(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L10D));
DFF_save_fm DFF_W3658(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L11D));
DFF_save_fm DFF_W3659(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L12D));
DFF_save_fm DFF_W3660(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L20D));
DFF_save_fm DFF_W3661(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L21D));
DFF_save_fm DFF_W3662(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L22D));
DFF_save_fm DFF_W3663(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L00E));
DFF_save_fm DFF_W3664(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L01E));
DFF_save_fm DFF_W3665(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L02E));
DFF_save_fm DFF_W3666(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L10E));
DFF_save_fm DFF_W3667(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L11E));
DFF_save_fm DFF_W3668(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L12E));
DFF_save_fm DFF_W3669(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L20E));
DFF_save_fm DFF_W3670(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L21E));
DFF_save_fm DFF_W3671(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L22E));
DFF_save_fm DFF_W3672(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L00F));
DFF_save_fm DFF_W3673(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L01F));
DFF_save_fm DFF_W3674(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2L02F));
DFF_save_fm DFF_W3675(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L10F));
DFF_save_fm DFF_W3676(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L11F));
DFF_save_fm DFF_W3677(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L12F));
DFF_save_fm DFF_W3678(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L20F));
DFF_save_fm DFF_W3679(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L21F));
DFF_save_fm DFF_W3680(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2L22F));
DFF_save_fm DFF_W3681(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M000));
DFF_save_fm DFF_W3682(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M010));
DFF_save_fm DFF_W3683(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M020));
DFF_save_fm DFF_W3684(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M100));
DFF_save_fm DFF_W3685(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M110));
DFF_save_fm DFF_W3686(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M120));
DFF_save_fm DFF_W3687(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M200));
DFF_save_fm DFF_W3688(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M210));
DFF_save_fm DFF_W3689(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M220));
DFF_save_fm DFF_W3690(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M001));
DFF_save_fm DFF_W3691(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M011));
DFF_save_fm DFF_W3692(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M021));
DFF_save_fm DFF_W3693(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M101));
DFF_save_fm DFF_W3694(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M111));
DFF_save_fm DFF_W3695(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M121));
DFF_save_fm DFF_W3696(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M201));
DFF_save_fm DFF_W3697(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M211));
DFF_save_fm DFF_W3698(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M221));
DFF_save_fm DFF_W3699(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M002));
DFF_save_fm DFF_W3700(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M012));
DFF_save_fm DFF_W3701(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M022));
DFF_save_fm DFF_W3702(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M102));
DFF_save_fm DFF_W3703(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M112));
DFF_save_fm DFF_W3704(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M122));
DFF_save_fm DFF_W3705(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M202));
DFF_save_fm DFF_W3706(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M212));
DFF_save_fm DFF_W3707(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M222));
DFF_save_fm DFF_W3708(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M003));
DFF_save_fm DFF_W3709(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M013));
DFF_save_fm DFF_W3710(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M023));
DFF_save_fm DFF_W3711(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M103));
DFF_save_fm DFF_W3712(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M113));
DFF_save_fm DFF_W3713(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M123));
DFF_save_fm DFF_W3714(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M203));
DFF_save_fm DFF_W3715(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M213));
DFF_save_fm DFF_W3716(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M223));
DFF_save_fm DFF_W3717(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M004));
DFF_save_fm DFF_W3718(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M014));
DFF_save_fm DFF_W3719(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M024));
DFF_save_fm DFF_W3720(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M104));
DFF_save_fm DFF_W3721(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M114));
DFF_save_fm DFF_W3722(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M124));
DFF_save_fm DFF_W3723(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M204));
DFF_save_fm DFF_W3724(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M214));
DFF_save_fm DFF_W3725(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M224));
DFF_save_fm DFF_W3726(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M005));
DFF_save_fm DFF_W3727(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M015));
DFF_save_fm DFF_W3728(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M025));
DFF_save_fm DFF_W3729(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M105));
DFF_save_fm DFF_W3730(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M115));
DFF_save_fm DFF_W3731(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M125));
DFF_save_fm DFF_W3732(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M205));
DFF_save_fm DFF_W3733(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M215));
DFF_save_fm DFF_W3734(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M225));
DFF_save_fm DFF_W3735(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M006));
DFF_save_fm DFF_W3736(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M016));
DFF_save_fm DFF_W3737(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M026));
DFF_save_fm DFF_W3738(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M106));
DFF_save_fm DFF_W3739(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M116));
DFF_save_fm DFF_W3740(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M126));
DFF_save_fm DFF_W3741(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M206));
DFF_save_fm DFF_W3742(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M216));
DFF_save_fm DFF_W3743(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M226));
DFF_save_fm DFF_W3744(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M007));
DFF_save_fm DFF_W3745(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M017));
DFF_save_fm DFF_W3746(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M027));
DFF_save_fm DFF_W3747(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M107));
DFF_save_fm DFF_W3748(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M117));
DFF_save_fm DFF_W3749(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M127));
DFF_save_fm DFF_W3750(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M207));
DFF_save_fm DFF_W3751(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M217));
DFF_save_fm DFF_W3752(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M227));
DFF_save_fm DFF_W3753(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M008));
DFF_save_fm DFF_W3754(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M018));
DFF_save_fm DFF_W3755(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M028));
DFF_save_fm DFF_W3756(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M108));
DFF_save_fm DFF_W3757(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M118));
DFF_save_fm DFF_W3758(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M128));
DFF_save_fm DFF_W3759(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M208));
DFF_save_fm DFF_W3760(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M218));
DFF_save_fm DFF_W3761(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M228));
DFF_save_fm DFF_W3762(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M009));
DFF_save_fm DFF_W3763(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M019));
DFF_save_fm DFF_W3764(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M029));
DFF_save_fm DFF_W3765(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M109));
DFF_save_fm DFF_W3766(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M119));
DFF_save_fm DFF_W3767(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M129));
DFF_save_fm DFF_W3768(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M209));
DFF_save_fm DFF_W3769(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M219));
DFF_save_fm DFF_W3770(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M229));
DFF_save_fm DFF_W3771(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M00A));
DFF_save_fm DFF_W3772(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M01A));
DFF_save_fm DFF_W3773(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M02A));
DFF_save_fm DFF_W3774(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M10A));
DFF_save_fm DFF_W3775(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M11A));
DFF_save_fm DFF_W3776(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M12A));
DFF_save_fm DFF_W3777(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M20A));
DFF_save_fm DFF_W3778(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M21A));
DFF_save_fm DFF_W3779(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M22A));
DFF_save_fm DFF_W3780(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M00B));
DFF_save_fm DFF_W3781(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M01B));
DFF_save_fm DFF_W3782(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M02B));
DFF_save_fm DFF_W3783(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M10B));
DFF_save_fm DFF_W3784(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M11B));
DFF_save_fm DFF_W3785(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M12B));
DFF_save_fm DFF_W3786(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M20B));
DFF_save_fm DFF_W3787(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M21B));
DFF_save_fm DFF_W3788(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M22B));
DFF_save_fm DFF_W3789(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M00C));
DFF_save_fm DFF_W3790(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M01C));
DFF_save_fm DFF_W3791(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M02C));
DFF_save_fm DFF_W3792(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M10C));
DFF_save_fm DFF_W3793(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M11C));
DFF_save_fm DFF_W3794(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M12C));
DFF_save_fm DFF_W3795(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M20C));
DFF_save_fm DFF_W3796(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M21C));
DFF_save_fm DFF_W3797(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M22C));
DFF_save_fm DFF_W3798(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M00D));
DFF_save_fm DFF_W3799(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M01D));
DFF_save_fm DFF_W3800(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M02D));
DFF_save_fm DFF_W3801(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M10D));
DFF_save_fm DFF_W3802(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M11D));
DFF_save_fm DFF_W3803(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M12D));
DFF_save_fm DFF_W3804(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M20D));
DFF_save_fm DFF_W3805(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M21D));
DFF_save_fm DFF_W3806(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M22D));
DFF_save_fm DFF_W3807(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M00E));
DFF_save_fm DFF_W3808(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M01E));
DFF_save_fm DFF_W3809(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M02E));
DFF_save_fm DFF_W3810(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M10E));
DFF_save_fm DFF_W3811(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M11E));
DFF_save_fm DFF_W3812(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M12E));
DFF_save_fm DFF_W3813(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M20E));
DFF_save_fm DFF_W3814(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M21E));
DFF_save_fm DFF_W3815(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M22E));
DFF_save_fm DFF_W3816(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M00F));
DFF_save_fm DFF_W3817(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M01F));
DFF_save_fm DFF_W3818(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M02F));
DFF_save_fm DFF_W3819(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M10F));
DFF_save_fm DFF_W3820(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2M11F));
DFF_save_fm DFF_W3821(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M12F));
DFF_save_fm DFF_W3822(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M20F));
DFF_save_fm DFF_W3823(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M21F));
DFF_save_fm DFF_W3824(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2M22F));
DFF_save_fm DFF_W3825(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N000));
DFF_save_fm DFF_W3826(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N010));
DFF_save_fm DFF_W3827(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N020));
DFF_save_fm DFF_W3828(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N100));
DFF_save_fm DFF_W3829(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N110));
DFF_save_fm DFF_W3830(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N120));
DFF_save_fm DFF_W3831(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N200));
DFF_save_fm DFF_W3832(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N210));
DFF_save_fm DFF_W3833(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N220));
DFF_save_fm DFF_W3834(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N001));
DFF_save_fm DFF_W3835(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N011));
DFF_save_fm DFF_W3836(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N021));
DFF_save_fm DFF_W3837(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N101));
DFF_save_fm DFF_W3838(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N111));
DFF_save_fm DFF_W3839(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N121));
DFF_save_fm DFF_W3840(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N201));
DFF_save_fm DFF_W3841(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N211));
DFF_save_fm DFF_W3842(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N221));
DFF_save_fm DFF_W3843(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N002));
DFF_save_fm DFF_W3844(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N012));
DFF_save_fm DFF_W3845(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N022));
DFF_save_fm DFF_W3846(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N102));
DFF_save_fm DFF_W3847(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N112));
DFF_save_fm DFF_W3848(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N122));
DFF_save_fm DFF_W3849(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N202));
DFF_save_fm DFF_W3850(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N212));
DFF_save_fm DFF_W3851(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N222));
DFF_save_fm DFF_W3852(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N003));
DFF_save_fm DFF_W3853(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N013));
DFF_save_fm DFF_W3854(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N023));
DFF_save_fm DFF_W3855(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N103));
DFF_save_fm DFF_W3856(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N113));
DFF_save_fm DFF_W3857(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N123));
DFF_save_fm DFF_W3858(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N203));
DFF_save_fm DFF_W3859(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N213));
DFF_save_fm DFF_W3860(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N223));
DFF_save_fm DFF_W3861(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N004));
DFF_save_fm DFF_W3862(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N014));
DFF_save_fm DFF_W3863(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N024));
DFF_save_fm DFF_W3864(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N104));
DFF_save_fm DFF_W3865(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N114));
DFF_save_fm DFF_W3866(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N124));
DFF_save_fm DFF_W3867(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N204));
DFF_save_fm DFF_W3868(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N214));
DFF_save_fm DFF_W3869(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N224));
DFF_save_fm DFF_W3870(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N005));
DFF_save_fm DFF_W3871(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N015));
DFF_save_fm DFF_W3872(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N025));
DFF_save_fm DFF_W3873(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N105));
DFF_save_fm DFF_W3874(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N115));
DFF_save_fm DFF_W3875(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N125));
DFF_save_fm DFF_W3876(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N205));
DFF_save_fm DFF_W3877(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N215));
DFF_save_fm DFF_W3878(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N225));
DFF_save_fm DFF_W3879(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N006));
DFF_save_fm DFF_W3880(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N016));
DFF_save_fm DFF_W3881(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N026));
DFF_save_fm DFF_W3882(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N106));
DFF_save_fm DFF_W3883(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N116));
DFF_save_fm DFF_W3884(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N126));
DFF_save_fm DFF_W3885(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N206));
DFF_save_fm DFF_W3886(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N216));
DFF_save_fm DFF_W3887(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N226));
DFF_save_fm DFF_W3888(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N007));
DFF_save_fm DFF_W3889(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N017));
DFF_save_fm DFF_W3890(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N027));
DFF_save_fm DFF_W3891(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N107));
DFF_save_fm DFF_W3892(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N117));
DFF_save_fm DFF_W3893(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N127));
DFF_save_fm DFF_W3894(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N207));
DFF_save_fm DFF_W3895(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N217));
DFF_save_fm DFF_W3896(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N227));
DFF_save_fm DFF_W3897(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N008));
DFF_save_fm DFF_W3898(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N018));
DFF_save_fm DFF_W3899(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N028));
DFF_save_fm DFF_W3900(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N108));
DFF_save_fm DFF_W3901(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N118));
DFF_save_fm DFF_W3902(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N128));
DFF_save_fm DFF_W3903(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N208));
DFF_save_fm DFF_W3904(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N218));
DFF_save_fm DFF_W3905(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N228));
DFF_save_fm DFF_W3906(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N009));
DFF_save_fm DFF_W3907(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N019));
DFF_save_fm DFF_W3908(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N029));
DFF_save_fm DFF_W3909(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N109));
DFF_save_fm DFF_W3910(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N119));
DFF_save_fm DFF_W3911(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N129));
DFF_save_fm DFF_W3912(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N209));
DFF_save_fm DFF_W3913(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N219));
DFF_save_fm DFF_W3914(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N229));
DFF_save_fm DFF_W3915(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N00A));
DFF_save_fm DFF_W3916(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N01A));
DFF_save_fm DFF_W3917(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N02A));
DFF_save_fm DFF_W3918(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N10A));
DFF_save_fm DFF_W3919(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N11A));
DFF_save_fm DFF_W3920(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N12A));
DFF_save_fm DFF_W3921(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N20A));
DFF_save_fm DFF_W3922(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N21A));
DFF_save_fm DFF_W3923(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N22A));
DFF_save_fm DFF_W3924(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N00B));
DFF_save_fm DFF_W3925(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N01B));
DFF_save_fm DFF_W3926(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N02B));
DFF_save_fm DFF_W3927(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N10B));
DFF_save_fm DFF_W3928(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N11B));
DFF_save_fm DFF_W3929(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N12B));
DFF_save_fm DFF_W3930(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N20B));
DFF_save_fm DFF_W3931(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N21B));
DFF_save_fm DFF_W3932(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N22B));
DFF_save_fm DFF_W3933(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N00C));
DFF_save_fm DFF_W3934(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N01C));
DFF_save_fm DFF_W3935(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N02C));
DFF_save_fm DFF_W3936(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N10C));
DFF_save_fm DFF_W3937(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N11C));
DFF_save_fm DFF_W3938(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N12C));
DFF_save_fm DFF_W3939(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N20C));
DFF_save_fm DFF_W3940(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N21C));
DFF_save_fm DFF_W3941(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N22C));
DFF_save_fm DFF_W3942(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N00D));
DFF_save_fm DFF_W3943(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N01D));
DFF_save_fm DFF_W3944(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N02D));
DFF_save_fm DFF_W3945(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N10D));
DFF_save_fm DFF_W3946(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N11D));
DFF_save_fm DFF_W3947(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N12D));
DFF_save_fm DFF_W3948(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N20D));
DFF_save_fm DFF_W3949(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N21D));
DFF_save_fm DFF_W3950(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N22D));
DFF_save_fm DFF_W3951(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N00E));
DFF_save_fm DFF_W3952(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N01E));
DFF_save_fm DFF_W3953(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N02E));
DFF_save_fm DFF_W3954(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N10E));
DFF_save_fm DFF_W3955(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N11E));
DFF_save_fm DFF_W3956(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N12E));
DFF_save_fm DFF_W3957(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N20E));
DFF_save_fm DFF_W3958(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N21E));
DFF_save_fm DFF_W3959(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N22E));
DFF_save_fm DFF_W3960(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N00F));
DFF_save_fm DFF_W3961(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N01F));
DFF_save_fm DFF_W3962(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N02F));
DFF_save_fm DFF_W3963(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N10F));
DFF_save_fm DFF_W3964(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N11F));
DFF_save_fm DFF_W3965(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N12F));
DFF_save_fm DFF_W3966(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N20F));
DFF_save_fm DFF_W3967(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2N21F));
DFF_save_fm DFF_W3968(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2N22F));
DFF_save_fm DFF_W3969(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O000));
DFF_save_fm DFF_W3970(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O010));
DFF_save_fm DFF_W3971(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O020));
DFF_save_fm DFF_W3972(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O100));
DFF_save_fm DFF_W3973(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O110));
DFF_save_fm DFF_W3974(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O120));
DFF_save_fm DFF_W3975(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O200));
DFF_save_fm DFF_W3976(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O210));
DFF_save_fm DFF_W3977(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O220));
DFF_save_fm DFF_W3978(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O001));
DFF_save_fm DFF_W3979(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O011));
DFF_save_fm DFF_W3980(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O021));
DFF_save_fm DFF_W3981(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O101));
DFF_save_fm DFF_W3982(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O111));
DFF_save_fm DFF_W3983(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O121));
DFF_save_fm DFF_W3984(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O201));
DFF_save_fm DFF_W3985(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O211));
DFF_save_fm DFF_W3986(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O221));
DFF_save_fm DFF_W3987(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O002));
DFF_save_fm DFF_W3988(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O012));
DFF_save_fm DFF_W3989(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O022));
DFF_save_fm DFF_W3990(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O102));
DFF_save_fm DFF_W3991(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O112));
DFF_save_fm DFF_W3992(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O122));
DFF_save_fm DFF_W3993(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O202));
DFF_save_fm DFF_W3994(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O212));
DFF_save_fm DFF_W3995(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O222));
DFF_save_fm DFF_W3996(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O003));
DFF_save_fm DFF_W3997(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O013));
DFF_save_fm DFF_W3998(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O023));
DFF_save_fm DFF_W3999(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O103));
DFF_save_fm DFF_W4000(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O113));
DFF_save_fm DFF_W4001(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O123));
DFF_save_fm DFF_W4002(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O203));
DFF_save_fm DFF_W4003(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O213));
DFF_save_fm DFF_W4004(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O223));
DFF_save_fm DFF_W4005(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O004));
DFF_save_fm DFF_W4006(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O014));
DFF_save_fm DFF_W4007(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O024));
DFF_save_fm DFF_W4008(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O104));
DFF_save_fm DFF_W4009(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O114));
DFF_save_fm DFF_W4010(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O124));
DFF_save_fm DFF_W4011(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O204));
DFF_save_fm DFF_W4012(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O214));
DFF_save_fm DFF_W4013(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O224));
DFF_save_fm DFF_W4014(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O005));
DFF_save_fm DFF_W4015(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O015));
DFF_save_fm DFF_W4016(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O025));
DFF_save_fm DFF_W4017(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O105));
DFF_save_fm DFF_W4018(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O115));
DFF_save_fm DFF_W4019(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O125));
DFF_save_fm DFF_W4020(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O205));
DFF_save_fm DFF_W4021(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O215));
DFF_save_fm DFF_W4022(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O225));
DFF_save_fm DFF_W4023(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O006));
DFF_save_fm DFF_W4024(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O016));
DFF_save_fm DFF_W4025(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O026));
DFF_save_fm DFF_W4026(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O106));
DFF_save_fm DFF_W4027(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O116));
DFF_save_fm DFF_W4028(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O126));
DFF_save_fm DFF_W4029(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O206));
DFF_save_fm DFF_W4030(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O216));
DFF_save_fm DFF_W4031(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O226));
DFF_save_fm DFF_W4032(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O007));
DFF_save_fm DFF_W4033(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O017));
DFF_save_fm DFF_W4034(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O027));
DFF_save_fm DFF_W4035(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O107));
DFF_save_fm DFF_W4036(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O117));
DFF_save_fm DFF_W4037(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O127));
DFF_save_fm DFF_W4038(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O207));
DFF_save_fm DFF_W4039(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O217));
DFF_save_fm DFF_W4040(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O227));
DFF_save_fm DFF_W4041(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O008));
DFF_save_fm DFF_W4042(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O018));
DFF_save_fm DFF_W4043(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O028));
DFF_save_fm DFF_W4044(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O108));
DFF_save_fm DFF_W4045(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O118));
DFF_save_fm DFF_W4046(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O128));
DFF_save_fm DFF_W4047(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O208));
DFF_save_fm DFF_W4048(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O218));
DFF_save_fm DFF_W4049(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O228));
DFF_save_fm DFF_W4050(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O009));
DFF_save_fm DFF_W4051(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O019));
DFF_save_fm DFF_W4052(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O029));
DFF_save_fm DFF_W4053(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O109));
DFF_save_fm DFF_W4054(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O119));
DFF_save_fm DFF_W4055(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O129));
DFF_save_fm DFF_W4056(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O209));
DFF_save_fm DFF_W4057(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O219));
DFF_save_fm DFF_W4058(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O229));
DFF_save_fm DFF_W4059(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O00A));
DFF_save_fm DFF_W4060(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O01A));
DFF_save_fm DFF_W4061(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O02A));
DFF_save_fm DFF_W4062(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O10A));
DFF_save_fm DFF_W4063(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O11A));
DFF_save_fm DFF_W4064(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O12A));
DFF_save_fm DFF_W4065(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O20A));
DFF_save_fm DFF_W4066(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O21A));
DFF_save_fm DFF_W4067(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O22A));
DFF_save_fm DFF_W4068(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O00B));
DFF_save_fm DFF_W4069(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O01B));
DFF_save_fm DFF_W4070(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O02B));
DFF_save_fm DFF_W4071(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O10B));
DFF_save_fm DFF_W4072(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O11B));
DFF_save_fm DFF_W4073(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O12B));
DFF_save_fm DFF_W4074(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O20B));
DFF_save_fm DFF_W4075(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O21B));
DFF_save_fm DFF_W4076(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O22B));
DFF_save_fm DFF_W4077(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O00C));
DFF_save_fm DFF_W4078(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O01C));
DFF_save_fm DFF_W4079(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O02C));
DFF_save_fm DFF_W4080(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O10C));
DFF_save_fm DFF_W4081(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O11C));
DFF_save_fm DFF_W4082(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O12C));
DFF_save_fm DFF_W4083(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O20C));
DFF_save_fm DFF_W4084(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O21C));
DFF_save_fm DFF_W4085(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O22C));
DFF_save_fm DFF_W4086(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O00D));
DFF_save_fm DFF_W4087(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O01D));
DFF_save_fm DFF_W4088(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O02D));
DFF_save_fm DFF_W4089(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O10D));
DFF_save_fm DFF_W4090(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O11D));
DFF_save_fm DFF_W4091(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O12D));
DFF_save_fm DFF_W4092(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O20D));
DFF_save_fm DFF_W4093(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O21D));
DFF_save_fm DFF_W4094(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O22D));
DFF_save_fm DFF_W4095(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O00E));
DFF_save_fm DFF_W4096(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O01E));
DFF_save_fm DFF_W4097(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O02E));
DFF_save_fm DFF_W4098(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O10E));
DFF_save_fm DFF_W4099(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O11E));
DFF_save_fm DFF_W4100(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O12E));
DFF_save_fm DFF_W4101(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O20E));
DFF_save_fm DFF_W4102(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O21E));
DFF_save_fm DFF_W4103(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O22E));
DFF_save_fm DFF_W4104(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O00F));
DFF_save_fm DFF_W4105(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O01F));
DFF_save_fm DFF_W4106(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O02F));
DFF_save_fm DFF_W4107(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O10F));
DFF_save_fm DFF_W4108(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O11F));
DFF_save_fm DFF_W4109(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2O12F));
DFF_save_fm DFF_W4110(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O20F));
DFF_save_fm DFF_W4111(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O21F));
DFF_save_fm DFF_W4112(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2O22F));
DFF_save_fm DFF_W4113(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P000));
DFF_save_fm DFF_W4114(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P010));
DFF_save_fm DFF_W4115(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P020));
DFF_save_fm DFF_W4116(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P100));
DFF_save_fm DFF_W4117(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P110));
DFF_save_fm DFF_W4118(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P120));
DFF_save_fm DFF_W4119(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P200));
DFF_save_fm DFF_W4120(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P210));
DFF_save_fm DFF_W4121(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P220));
DFF_save_fm DFF_W4122(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P001));
DFF_save_fm DFF_W4123(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P011));
DFF_save_fm DFF_W4124(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P021));
DFF_save_fm DFF_W4125(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P101));
DFF_save_fm DFF_W4126(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P111));
DFF_save_fm DFF_W4127(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P121));
DFF_save_fm DFF_W4128(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P201));
DFF_save_fm DFF_W4129(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P211));
DFF_save_fm DFF_W4130(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P221));
DFF_save_fm DFF_W4131(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P002));
DFF_save_fm DFF_W4132(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P012));
DFF_save_fm DFF_W4133(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P022));
DFF_save_fm DFF_W4134(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P102));
DFF_save_fm DFF_W4135(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P112));
DFF_save_fm DFF_W4136(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P122));
DFF_save_fm DFF_W4137(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P202));
DFF_save_fm DFF_W4138(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P212));
DFF_save_fm DFF_W4139(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P222));
DFF_save_fm DFF_W4140(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P003));
DFF_save_fm DFF_W4141(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P013));
DFF_save_fm DFF_W4142(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P023));
DFF_save_fm DFF_W4143(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P103));
DFF_save_fm DFF_W4144(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P113));
DFF_save_fm DFF_W4145(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P123));
DFF_save_fm DFF_W4146(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P203));
DFF_save_fm DFF_W4147(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P213));
DFF_save_fm DFF_W4148(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P223));
DFF_save_fm DFF_W4149(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P004));
DFF_save_fm DFF_W4150(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P014));
DFF_save_fm DFF_W4151(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P024));
DFF_save_fm DFF_W4152(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P104));
DFF_save_fm DFF_W4153(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P114));
DFF_save_fm DFF_W4154(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P124));
DFF_save_fm DFF_W4155(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P204));
DFF_save_fm DFF_W4156(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P214));
DFF_save_fm DFF_W4157(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P224));
DFF_save_fm DFF_W4158(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P005));
DFF_save_fm DFF_W4159(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P015));
DFF_save_fm DFF_W4160(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P025));
DFF_save_fm DFF_W4161(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P105));
DFF_save_fm DFF_W4162(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P115));
DFF_save_fm DFF_W4163(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P125));
DFF_save_fm DFF_W4164(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P205));
DFF_save_fm DFF_W4165(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P215));
DFF_save_fm DFF_W4166(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P225));
DFF_save_fm DFF_W4167(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P006));
DFF_save_fm DFF_W4168(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P016));
DFF_save_fm DFF_W4169(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P026));
DFF_save_fm DFF_W4170(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P106));
DFF_save_fm DFF_W4171(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P116));
DFF_save_fm DFF_W4172(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P126));
DFF_save_fm DFF_W4173(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P206));
DFF_save_fm DFF_W4174(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P216));
DFF_save_fm DFF_W4175(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P226));
DFF_save_fm DFF_W4176(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P007));
DFF_save_fm DFF_W4177(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P017));
DFF_save_fm DFF_W4178(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P027));
DFF_save_fm DFF_W4179(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P107));
DFF_save_fm DFF_W4180(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P117));
DFF_save_fm DFF_W4181(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P127));
DFF_save_fm DFF_W4182(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P207));
DFF_save_fm DFF_W4183(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P217));
DFF_save_fm DFF_W4184(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P227));
DFF_save_fm DFF_W4185(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P008));
DFF_save_fm DFF_W4186(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P018));
DFF_save_fm DFF_W4187(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P028));
DFF_save_fm DFF_W4188(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P108));
DFF_save_fm DFF_W4189(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P118));
DFF_save_fm DFF_W4190(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P128));
DFF_save_fm DFF_W4191(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P208));
DFF_save_fm DFF_W4192(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P218));
DFF_save_fm DFF_W4193(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P228));
DFF_save_fm DFF_W4194(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P009));
DFF_save_fm DFF_W4195(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P019));
DFF_save_fm DFF_W4196(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P029));
DFF_save_fm DFF_W4197(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P109));
DFF_save_fm DFF_W4198(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P119));
DFF_save_fm DFF_W4199(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P129));
DFF_save_fm DFF_W4200(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P209));
DFF_save_fm DFF_W4201(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P219));
DFF_save_fm DFF_W4202(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P229));
DFF_save_fm DFF_W4203(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P00A));
DFF_save_fm DFF_W4204(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P01A));
DFF_save_fm DFF_W4205(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P02A));
DFF_save_fm DFF_W4206(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P10A));
DFF_save_fm DFF_W4207(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P11A));
DFF_save_fm DFF_W4208(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P12A));
DFF_save_fm DFF_W4209(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P20A));
DFF_save_fm DFF_W4210(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P21A));
DFF_save_fm DFF_W4211(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P22A));
DFF_save_fm DFF_W4212(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P00B));
DFF_save_fm DFF_W4213(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P01B));
DFF_save_fm DFF_W4214(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P02B));
DFF_save_fm DFF_W4215(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P10B));
DFF_save_fm DFF_W4216(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P11B));
DFF_save_fm DFF_W4217(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P12B));
DFF_save_fm DFF_W4218(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P20B));
DFF_save_fm DFF_W4219(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P21B));
DFF_save_fm DFF_W4220(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P22B));
DFF_save_fm DFF_W4221(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P00C));
DFF_save_fm DFF_W4222(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P01C));
DFF_save_fm DFF_W4223(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P02C));
DFF_save_fm DFF_W4224(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P10C));
DFF_save_fm DFF_W4225(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P11C));
DFF_save_fm DFF_W4226(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P12C));
DFF_save_fm DFF_W4227(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P20C));
DFF_save_fm DFF_W4228(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P21C));
DFF_save_fm DFF_W4229(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P22C));
DFF_save_fm DFF_W4230(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P00D));
DFF_save_fm DFF_W4231(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P01D));
DFF_save_fm DFF_W4232(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P02D));
DFF_save_fm DFF_W4233(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P10D));
DFF_save_fm DFF_W4234(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P11D));
DFF_save_fm DFF_W4235(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P12D));
DFF_save_fm DFF_W4236(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P20D));
DFF_save_fm DFF_W4237(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P21D));
DFF_save_fm DFF_W4238(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P22D));
DFF_save_fm DFF_W4239(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P00E));
DFF_save_fm DFF_W4240(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P01E));
DFF_save_fm DFF_W4241(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P02E));
DFF_save_fm DFF_W4242(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P10E));
DFF_save_fm DFF_W4243(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P11E));
DFF_save_fm DFF_W4244(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P12E));
DFF_save_fm DFF_W4245(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P20E));
DFF_save_fm DFF_W4246(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P21E));
DFF_save_fm DFF_W4247(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P22E));
DFF_save_fm DFF_W4248(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P00F));
DFF_save_fm DFF_W4249(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P01F));
DFF_save_fm DFF_W4250(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P02F));
DFF_save_fm DFF_W4251(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P10F));
DFF_save_fm DFF_W4252(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P11F));
DFF_save_fm DFF_W4253(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P12F));
DFF_save_fm DFF_W4254(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2P20F));
DFF_save_fm DFF_W4255(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P21F));
DFF_save_fm DFF_W4256(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2P22F));
DFF_save_fm DFF_W4257(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q000));
DFF_save_fm DFF_W4258(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q010));
DFF_save_fm DFF_W4259(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q020));
DFF_save_fm DFF_W4260(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q100));
DFF_save_fm DFF_W4261(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q110));
DFF_save_fm DFF_W4262(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q120));
DFF_save_fm DFF_W4263(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q200));
DFF_save_fm DFF_W4264(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q210));
DFF_save_fm DFF_W4265(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q220));
DFF_save_fm DFF_W4266(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q001));
DFF_save_fm DFF_W4267(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q011));
DFF_save_fm DFF_W4268(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q021));
DFF_save_fm DFF_W4269(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q101));
DFF_save_fm DFF_W4270(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q111));
DFF_save_fm DFF_W4271(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q121));
DFF_save_fm DFF_W4272(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q201));
DFF_save_fm DFF_W4273(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q211));
DFF_save_fm DFF_W4274(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q221));
DFF_save_fm DFF_W4275(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q002));
DFF_save_fm DFF_W4276(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q012));
DFF_save_fm DFF_W4277(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q022));
DFF_save_fm DFF_W4278(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q102));
DFF_save_fm DFF_W4279(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q112));
DFF_save_fm DFF_W4280(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q122));
DFF_save_fm DFF_W4281(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q202));
DFF_save_fm DFF_W4282(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q212));
DFF_save_fm DFF_W4283(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q222));
DFF_save_fm DFF_W4284(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q003));
DFF_save_fm DFF_W4285(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q013));
DFF_save_fm DFF_W4286(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q023));
DFF_save_fm DFF_W4287(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q103));
DFF_save_fm DFF_W4288(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q113));
DFF_save_fm DFF_W4289(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q123));
DFF_save_fm DFF_W4290(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q203));
DFF_save_fm DFF_W4291(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q213));
DFF_save_fm DFF_W4292(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q223));
DFF_save_fm DFF_W4293(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q004));
DFF_save_fm DFF_W4294(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q014));
DFF_save_fm DFF_W4295(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q024));
DFF_save_fm DFF_W4296(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q104));
DFF_save_fm DFF_W4297(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q114));
DFF_save_fm DFF_W4298(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q124));
DFF_save_fm DFF_W4299(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q204));
DFF_save_fm DFF_W4300(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q214));
DFF_save_fm DFF_W4301(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q224));
DFF_save_fm DFF_W4302(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q005));
DFF_save_fm DFF_W4303(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q015));
DFF_save_fm DFF_W4304(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q025));
DFF_save_fm DFF_W4305(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q105));
DFF_save_fm DFF_W4306(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q115));
DFF_save_fm DFF_W4307(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q125));
DFF_save_fm DFF_W4308(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q205));
DFF_save_fm DFF_W4309(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q215));
DFF_save_fm DFF_W4310(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q225));
DFF_save_fm DFF_W4311(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q006));
DFF_save_fm DFF_W4312(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q016));
DFF_save_fm DFF_W4313(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q026));
DFF_save_fm DFF_W4314(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q106));
DFF_save_fm DFF_W4315(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q116));
DFF_save_fm DFF_W4316(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q126));
DFF_save_fm DFF_W4317(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q206));
DFF_save_fm DFF_W4318(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q216));
DFF_save_fm DFF_W4319(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q226));
DFF_save_fm DFF_W4320(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q007));
DFF_save_fm DFF_W4321(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q017));
DFF_save_fm DFF_W4322(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q027));
DFF_save_fm DFF_W4323(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q107));
DFF_save_fm DFF_W4324(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q117));
DFF_save_fm DFF_W4325(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q127));
DFF_save_fm DFF_W4326(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q207));
DFF_save_fm DFF_W4327(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q217));
DFF_save_fm DFF_W4328(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q227));
DFF_save_fm DFF_W4329(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q008));
DFF_save_fm DFF_W4330(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q018));
DFF_save_fm DFF_W4331(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q028));
DFF_save_fm DFF_W4332(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q108));
DFF_save_fm DFF_W4333(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q118));
DFF_save_fm DFF_W4334(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q128));
DFF_save_fm DFF_W4335(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q208));
DFF_save_fm DFF_W4336(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q218));
DFF_save_fm DFF_W4337(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q228));
DFF_save_fm DFF_W4338(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q009));
DFF_save_fm DFF_W4339(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q019));
DFF_save_fm DFF_W4340(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q029));
DFF_save_fm DFF_W4341(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q109));
DFF_save_fm DFF_W4342(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q119));
DFF_save_fm DFF_W4343(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q129));
DFF_save_fm DFF_W4344(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q209));
DFF_save_fm DFF_W4345(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q219));
DFF_save_fm DFF_W4346(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q229));
DFF_save_fm DFF_W4347(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q00A));
DFF_save_fm DFF_W4348(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q01A));
DFF_save_fm DFF_W4349(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q02A));
DFF_save_fm DFF_W4350(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q10A));
DFF_save_fm DFF_W4351(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q11A));
DFF_save_fm DFF_W4352(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q12A));
DFF_save_fm DFF_W4353(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q20A));
DFF_save_fm DFF_W4354(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q21A));
DFF_save_fm DFF_W4355(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q22A));
DFF_save_fm DFF_W4356(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q00B));
DFF_save_fm DFF_W4357(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q01B));
DFF_save_fm DFF_W4358(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q02B));
DFF_save_fm DFF_W4359(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q10B));
DFF_save_fm DFF_W4360(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q11B));
DFF_save_fm DFF_W4361(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q12B));
DFF_save_fm DFF_W4362(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q20B));
DFF_save_fm DFF_W4363(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q21B));
DFF_save_fm DFF_W4364(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q22B));
DFF_save_fm DFF_W4365(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q00C));
DFF_save_fm DFF_W4366(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q01C));
DFF_save_fm DFF_W4367(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q02C));
DFF_save_fm DFF_W4368(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q10C));
DFF_save_fm DFF_W4369(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q11C));
DFF_save_fm DFF_W4370(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q12C));
DFF_save_fm DFF_W4371(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q20C));
DFF_save_fm DFF_W4372(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q21C));
DFF_save_fm DFF_W4373(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q22C));
DFF_save_fm DFF_W4374(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q00D));
DFF_save_fm DFF_W4375(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q01D));
DFF_save_fm DFF_W4376(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q02D));
DFF_save_fm DFF_W4377(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q10D));
DFF_save_fm DFF_W4378(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q11D));
DFF_save_fm DFF_W4379(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q12D));
DFF_save_fm DFF_W4380(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q20D));
DFF_save_fm DFF_W4381(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q21D));
DFF_save_fm DFF_W4382(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q22D));
DFF_save_fm DFF_W4383(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q00E));
DFF_save_fm DFF_W4384(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q01E));
DFF_save_fm DFF_W4385(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q02E));
DFF_save_fm DFF_W4386(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q10E));
DFF_save_fm DFF_W4387(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q11E));
DFF_save_fm DFF_W4388(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q12E));
DFF_save_fm DFF_W4389(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q20E));
DFF_save_fm DFF_W4390(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q21E));
DFF_save_fm DFF_W4391(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q22E));
DFF_save_fm DFF_W4392(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q00F));
DFF_save_fm DFF_W4393(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q01F));
DFF_save_fm DFF_W4394(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q02F));
DFF_save_fm DFF_W4395(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q10F));
DFF_save_fm DFF_W4396(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q11F));
DFF_save_fm DFF_W4397(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q12F));
DFF_save_fm DFF_W4398(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q20F));
DFF_save_fm DFF_W4399(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2Q21F));
DFF_save_fm DFF_W4400(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2Q22F));
DFF_save_fm DFF_W4401(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R000));
DFF_save_fm DFF_W4402(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R010));
DFF_save_fm DFF_W4403(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R020));
DFF_save_fm DFF_W4404(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R100));
DFF_save_fm DFF_W4405(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R110));
DFF_save_fm DFF_W4406(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R120));
DFF_save_fm DFF_W4407(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R200));
DFF_save_fm DFF_W4408(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R210));
DFF_save_fm DFF_W4409(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R220));
DFF_save_fm DFF_W4410(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R001));
DFF_save_fm DFF_W4411(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R011));
DFF_save_fm DFF_W4412(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R021));
DFF_save_fm DFF_W4413(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R101));
DFF_save_fm DFF_W4414(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R111));
DFF_save_fm DFF_W4415(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R121));
DFF_save_fm DFF_W4416(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R201));
DFF_save_fm DFF_W4417(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R211));
DFF_save_fm DFF_W4418(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R221));
DFF_save_fm DFF_W4419(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R002));
DFF_save_fm DFF_W4420(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R012));
DFF_save_fm DFF_W4421(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R022));
DFF_save_fm DFF_W4422(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R102));
DFF_save_fm DFF_W4423(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R112));
DFF_save_fm DFF_W4424(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R122));
DFF_save_fm DFF_W4425(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R202));
DFF_save_fm DFF_W4426(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R212));
DFF_save_fm DFF_W4427(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R222));
DFF_save_fm DFF_W4428(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R003));
DFF_save_fm DFF_W4429(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R013));
DFF_save_fm DFF_W4430(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R023));
DFF_save_fm DFF_W4431(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R103));
DFF_save_fm DFF_W4432(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R113));
DFF_save_fm DFF_W4433(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R123));
DFF_save_fm DFF_W4434(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R203));
DFF_save_fm DFF_W4435(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R213));
DFF_save_fm DFF_W4436(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R223));
DFF_save_fm DFF_W4437(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R004));
DFF_save_fm DFF_W4438(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R014));
DFF_save_fm DFF_W4439(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R024));
DFF_save_fm DFF_W4440(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R104));
DFF_save_fm DFF_W4441(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R114));
DFF_save_fm DFF_W4442(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R124));
DFF_save_fm DFF_W4443(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R204));
DFF_save_fm DFF_W4444(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R214));
DFF_save_fm DFF_W4445(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R224));
DFF_save_fm DFF_W4446(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R005));
DFF_save_fm DFF_W4447(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R015));
DFF_save_fm DFF_W4448(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R025));
DFF_save_fm DFF_W4449(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R105));
DFF_save_fm DFF_W4450(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R115));
DFF_save_fm DFF_W4451(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R125));
DFF_save_fm DFF_W4452(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R205));
DFF_save_fm DFF_W4453(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R215));
DFF_save_fm DFF_W4454(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R225));
DFF_save_fm DFF_W4455(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R006));
DFF_save_fm DFF_W4456(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R016));
DFF_save_fm DFF_W4457(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R026));
DFF_save_fm DFF_W4458(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R106));
DFF_save_fm DFF_W4459(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R116));
DFF_save_fm DFF_W4460(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R126));
DFF_save_fm DFF_W4461(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R206));
DFF_save_fm DFF_W4462(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R216));
DFF_save_fm DFF_W4463(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R226));
DFF_save_fm DFF_W4464(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R007));
DFF_save_fm DFF_W4465(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R017));
DFF_save_fm DFF_W4466(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R027));
DFF_save_fm DFF_W4467(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R107));
DFF_save_fm DFF_W4468(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R117));
DFF_save_fm DFF_W4469(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R127));
DFF_save_fm DFF_W4470(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R207));
DFF_save_fm DFF_W4471(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R217));
DFF_save_fm DFF_W4472(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R227));
DFF_save_fm DFF_W4473(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R008));
DFF_save_fm DFF_W4474(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R018));
DFF_save_fm DFF_W4475(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R028));
DFF_save_fm DFF_W4476(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R108));
DFF_save_fm DFF_W4477(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R118));
DFF_save_fm DFF_W4478(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R128));
DFF_save_fm DFF_W4479(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R208));
DFF_save_fm DFF_W4480(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R218));
DFF_save_fm DFF_W4481(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R228));
DFF_save_fm DFF_W4482(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R009));
DFF_save_fm DFF_W4483(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R019));
DFF_save_fm DFF_W4484(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R029));
DFF_save_fm DFF_W4485(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R109));
DFF_save_fm DFF_W4486(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R119));
DFF_save_fm DFF_W4487(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R129));
DFF_save_fm DFF_W4488(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R209));
DFF_save_fm DFF_W4489(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R219));
DFF_save_fm DFF_W4490(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R229));
DFF_save_fm DFF_W4491(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R00A));
DFF_save_fm DFF_W4492(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R01A));
DFF_save_fm DFF_W4493(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R02A));
DFF_save_fm DFF_W4494(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R10A));
DFF_save_fm DFF_W4495(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R11A));
DFF_save_fm DFF_W4496(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R12A));
DFF_save_fm DFF_W4497(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R20A));
DFF_save_fm DFF_W4498(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R21A));
DFF_save_fm DFF_W4499(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R22A));
DFF_save_fm DFF_W4500(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R00B));
DFF_save_fm DFF_W4501(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R01B));
DFF_save_fm DFF_W4502(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R02B));
DFF_save_fm DFF_W4503(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R10B));
DFF_save_fm DFF_W4504(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R11B));
DFF_save_fm DFF_W4505(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R12B));
DFF_save_fm DFF_W4506(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R20B));
DFF_save_fm DFF_W4507(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R21B));
DFF_save_fm DFF_W4508(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R22B));
DFF_save_fm DFF_W4509(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R00C));
DFF_save_fm DFF_W4510(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R01C));
DFF_save_fm DFF_W4511(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R02C));
DFF_save_fm DFF_W4512(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R10C));
DFF_save_fm DFF_W4513(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R11C));
DFF_save_fm DFF_W4514(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R12C));
DFF_save_fm DFF_W4515(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R20C));
DFF_save_fm DFF_W4516(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R21C));
DFF_save_fm DFF_W4517(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R22C));
DFF_save_fm DFF_W4518(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R00D));
DFF_save_fm DFF_W4519(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R01D));
DFF_save_fm DFF_W4520(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R02D));
DFF_save_fm DFF_W4521(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R10D));
DFF_save_fm DFF_W4522(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R11D));
DFF_save_fm DFF_W4523(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R12D));
DFF_save_fm DFF_W4524(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R20D));
DFF_save_fm DFF_W4525(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R21D));
DFF_save_fm DFF_W4526(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R22D));
DFF_save_fm DFF_W4527(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R00E));
DFF_save_fm DFF_W4528(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R01E));
DFF_save_fm DFF_W4529(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R02E));
DFF_save_fm DFF_W4530(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R10E));
DFF_save_fm DFF_W4531(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R11E));
DFF_save_fm DFF_W4532(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R12E));
DFF_save_fm DFF_W4533(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R20E));
DFF_save_fm DFF_W4534(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R21E));
DFF_save_fm DFF_W4535(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R22E));
DFF_save_fm DFF_W4536(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R00F));
DFF_save_fm DFF_W4537(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R01F));
DFF_save_fm DFF_W4538(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R02F));
DFF_save_fm DFF_W4539(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R10F));
DFF_save_fm DFF_W4540(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R11F));
DFF_save_fm DFF_W4541(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2R12F));
DFF_save_fm DFF_W4542(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R20F));
DFF_save_fm DFF_W4543(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R21F));
DFF_save_fm DFF_W4544(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2R22F));
DFF_save_fm DFF_W4545(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S000));
DFF_save_fm DFF_W4546(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S010));
DFF_save_fm DFF_W4547(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S020));
DFF_save_fm DFF_W4548(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S100));
DFF_save_fm DFF_W4549(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S110));
DFF_save_fm DFF_W4550(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S120));
DFF_save_fm DFF_W4551(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S200));
DFF_save_fm DFF_W4552(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S210));
DFF_save_fm DFF_W4553(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S220));
DFF_save_fm DFF_W4554(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S001));
DFF_save_fm DFF_W4555(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S011));
DFF_save_fm DFF_W4556(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S021));
DFF_save_fm DFF_W4557(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S101));
DFF_save_fm DFF_W4558(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S111));
DFF_save_fm DFF_W4559(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S121));
DFF_save_fm DFF_W4560(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S201));
DFF_save_fm DFF_W4561(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S211));
DFF_save_fm DFF_W4562(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S221));
DFF_save_fm DFF_W4563(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S002));
DFF_save_fm DFF_W4564(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S012));
DFF_save_fm DFF_W4565(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S022));
DFF_save_fm DFF_W4566(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S102));
DFF_save_fm DFF_W4567(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S112));
DFF_save_fm DFF_W4568(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S122));
DFF_save_fm DFF_W4569(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S202));
DFF_save_fm DFF_W4570(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S212));
DFF_save_fm DFF_W4571(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S222));
DFF_save_fm DFF_W4572(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S003));
DFF_save_fm DFF_W4573(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S013));
DFF_save_fm DFF_W4574(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S023));
DFF_save_fm DFF_W4575(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S103));
DFF_save_fm DFF_W4576(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S113));
DFF_save_fm DFF_W4577(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S123));
DFF_save_fm DFF_W4578(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S203));
DFF_save_fm DFF_W4579(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S213));
DFF_save_fm DFF_W4580(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S223));
DFF_save_fm DFF_W4581(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S004));
DFF_save_fm DFF_W4582(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S014));
DFF_save_fm DFF_W4583(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S024));
DFF_save_fm DFF_W4584(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S104));
DFF_save_fm DFF_W4585(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S114));
DFF_save_fm DFF_W4586(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S124));
DFF_save_fm DFF_W4587(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S204));
DFF_save_fm DFF_W4588(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S214));
DFF_save_fm DFF_W4589(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S224));
DFF_save_fm DFF_W4590(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S005));
DFF_save_fm DFF_W4591(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S015));
DFF_save_fm DFF_W4592(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S025));
DFF_save_fm DFF_W4593(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S105));
DFF_save_fm DFF_W4594(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S115));
DFF_save_fm DFF_W4595(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S125));
DFF_save_fm DFF_W4596(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S205));
DFF_save_fm DFF_W4597(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S215));
DFF_save_fm DFF_W4598(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S225));
DFF_save_fm DFF_W4599(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S006));
DFF_save_fm DFF_W4600(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S016));
DFF_save_fm DFF_W4601(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S026));
DFF_save_fm DFF_W4602(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S106));
DFF_save_fm DFF_W4603(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S116));
DFF_save_fm DFF_W4604(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S126));
DFF_save_fm DFF_W4605(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S206));
DFF_save_fm DFF_W4606(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S216));
DFF_save_fm DFF_W4607(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S226));
DFF_save_fm DFF_W4608(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S007));
DFF_save_fm DFF_W4609(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S017));
DFF_save_fm DFF_W4610(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S027));
DFF_save_fm DFF_W4611(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S107));
DFF_save_fm DFF_W4612(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S117));
DFF_save_fm DFF_W4613(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S127));
DFF_save_fm DFF_W4614(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S207));
DFF_save_fm DFF_W4615(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S217));
DFF_save_fm DFF_W4616(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S227));
DFF_save_fm DFF_W4617(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S008));
DFF_save_fm DFF_W4618(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S018));
DFF_save_fm DFF_W4619(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S028));
DFF_save_fm DFF_W4620(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S108));
DFF_save_fm DFF_W4621(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S118));
DFF_save_fm DFF_W4622(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S128));
DFF_save_fm DFF_W4623(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S208));
DFF_save_fm DFF_W4624(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S218));
DFF_save_fm DFF_W4625(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S228));
DFF_save_fm DFF_W4626(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S009));
DFF_save_fm DFF_W4627(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S019));
DFF_save_fm DFF_W4628(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S029));
DFF_save_fm DFF_W4629(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S109));
DFF_save_fm DFF_W4630(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S119));
DFF_save_fm DFF_W4631(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S129));
DFF_save_fm DFF_W4632(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S209));
DFF_save_fm DFF_W4633(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S219));
DFF_save_fm DFF_W4634(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S229));
DFF_save_fm DFF_W4635(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S00A));
DFF_save_fm DFF_W4636(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S01A));
DFF_save_fm DFF_W4637(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S02A));
DFF_save_fm DFF_W4638(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S10A));
DFF_save_fm DFF_W4639(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S11A));
DFF_save_fm DFF_W4640(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S12A));
DFF_save_fm DFF_W4641(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S20A));
DFF_save_fm DFF_W4642(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S21A));
DFF_save_fm DFF_W4643(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S22A));
DFF_save_fm DFF_W4644(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S00B));
DFF_save_fm DFF_W4645(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S01B));
DFF_save_fm DFF_W4646(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S02B));
DFF_save_fm DFF_W4647(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S10B));
DFF_save_fm DFF_W4648(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S11B));
DFF_save_fm DFF_W4649(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S12B));
DFF_save_fm DFF_W4650(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S20B));
DFF_save_fm DFF_W4651(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S21B));
DFF_save_fm DFF_W4652(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S22B));
DFF_save_fm DFF_W4653(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S00C));
DFF_save_fm DFF_W4654(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S01C));
DFF_save_fm DFF_W4655(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S02C));
DFF_save_fm DFF_W4656(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S10C));
DFF_save_fm DFF_W4657(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S11C));
DFF_save_fm DFF_W4658(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S12C));
DFF_save_fm DFF_W4659(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S20C));
DFF_save_fm DFF_W4660(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S21C));
DFF_save_fm DFF_W4661(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S22C));
DFF_save_fm DFF_W4662(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S00D));
DFF_save_fm DFF_W4663(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S01D));
DFF_save_fm DFF_W4664(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S02D));
DFF_save_fm DFF_W4665(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S10D));
DFF_save_fm DFF_W4666(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S11D));
DFF_save_fm DFF_W4667(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S12D));
DFF_save_fm DFF_W4668(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S20D));
DFF_save_fm DFF_W4669(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S21D));
DFF_save_fm DFF_W4670(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S22D));
DFF_save_fm DFF_W4671(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S00E));
DFF_save_fm DFF_W4672(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S01E));
DFF_save_fm DFF_W4673(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S02E));
DFF_save_fm DFF_W4674(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S10E));
DFF_save_fm DFF_W4675(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S11E));
DFF_save_fm DFF_W4676(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S12E));
DFF_save_fm DFF_W4677(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S20E));
DFF_save_fm DFF_W4678(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S21E));
DFF_save_fm DFF_W4679(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S22E));
DFF_save_fm DFF_W4680(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S00F));
DFF_save_fm DFF_W4681(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S01F));
DFF_save_fm DFF_W4682(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S02F));
DFF_save_fm DFF_W4683(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S10F));
DFF_save_fm DFF_W4684(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S11F));
DFF_save_fm DFF_W4685(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S12F));
DFF_save_fm DFF_W4686(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S20F));
DFF_save_fm DFF_W4687(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2S21F));
DFF_save_fm DFF_W4688(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2S22F));
DFF_save_fm DFF_W4689(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T000));
DFF_save_fm DFF_W4690(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T010));
DFF_save_fm DFF_W4691(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T020));
DFF_save_fm DFF_W4692(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T100));
DFF_save_fm DFF_W4693(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T110));
DFF_save_fm DFF_W4694(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T120));
DFF_save_fm DFF_W4695(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T200));
DFF_save_fm DFF_W4696(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T210));
DFF_save_fm DFF_W4697(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T220));
DFF_save_fm DFF_W4698(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T001));
DFF_save_fm DFF_W4699(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T011));
DFF_save_fm DFF_W4700(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T021));
DFF_save_fm DFF_W4701(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T101));
DFF_save_fm DFF_W4702(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T111));
DFF_save_fm DFF_W4703(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T121));
DFF_save_fm DFF_W4704(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T201));
DFF_save_fm DFF_W4705(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T211));
DFF_save_fm DFF_W4706(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T221));
DFF_save_fm DFF_W4707(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T002));
DFF_save_fm DFF_W4708(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T012));
DFF_save_fm DFF_W4709(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T022));
DFF_save_fm DFF_W4710(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T102));
DFF_save_fm DFF_W4711(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T112));
DFF_save_fm DFF_W4712(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T122));
DFF_save_fm DFF_W4713(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T202));
DFF_save_fm DFF_W4714(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T212));
DFF_save_fm DFF_W4715(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T222));
DFF_save_fm DFF_W4716(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T003));
DFF_save_fm DFF_W4717(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T013));
DFF_save_fm DFF_W4718(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T023));
DFF_save_fm DFF_W4719(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T103));
DFF_save_fm DFF_W4720(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T113));
DFF_save_fm DFF_W4721(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T123));
DFF_save_fm DFF_W4722(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T203));
DFF_save_fm DFF_W4723(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T213));
DFF_save_fm DFF_W4724(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T223));
DFF_save_fm DFF_W4725(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T004));
DFF_save_fm DFF_W4726(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T014));
DFF_save_fm DFF_W4727(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T024));
DFF_save_fm DFF_W4728(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T104));
DFF_save_fm DFF_W4729(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T114));
DFF_save_fm DFF_W4730(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T124));
DFF_save_fm DFF_W4731(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T204));
DFF_save_fm DFF_W4732(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T214));
DFF_save_fm DFF_W4733(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T224));
DFF_save_fm DFF_W4734(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T005));
DFF_save_fm DFF_W4735(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T015));
DFF_save_fm DFF_W4736(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T025));
DFF_save_fm DFF_W4737(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T105));
DFF_save_fm DFF_W4738(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T115));
DFF_save_fm DFF_W4739(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T125));
DFF_save_fm DFF_W4740(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T205));
DFF_save_fm DFF_W4741(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T215));
DFF_save_fm DFF_W4742(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T225));
DFF_save_fm DFF_W4743(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T006));
DFF_save_fm DFF_W4744(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T016));
DFF_save_fm DFF_W4745(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T026));
DFF_save_fm DFF_W4746(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T106));
DFF_save_fm DFF_W4747(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T116));
DFF_save_fm DFF_W4748(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T126));
DFF_save_fm DFF_W4749(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T206));
DFF_save_fm DFF_W4750(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T216));
DFF_save_fm DFF_W4751(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T226));
DFF_save_fm DFF_W4752(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T007));
DFF_save_fm DFF_W4753(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T017));
DFF_save_fm DFF_W4754(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T027));
DFF_save_fm DFF_W4755(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T107));
DFF_save_fm DFF_W4756(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T117));
DFF_save_fm DFF_W4757(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T127));
DFF_save_fm DFF_W4758(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T207));
DFF_save_fm DFF_W4759(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T217));
DFF_save_fm DFF_W4760(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T227));
DFF_save_fm DFF_W4761(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T008));
DFF_save_fm DFF_W4762(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T018));
DFF_save_fm DFF_W4763(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T028));
DFF_save_fm DFF_W4764(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T108));
DFF_save_fm DFF_W4765(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T118));
DFF_save_fm DFF_W4766(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T128));
DFF_save_fm DFF_W4767(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T208));
DFF_save_fm DFF_W4768(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T218));
DFF_save_fm DFF_W4769(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T228));
DFF_save_fm DFF_W4770(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T009));
DFF_save_fm DFF_W4771(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T019));
DFF_save_fm DFF_W4772(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T029));
DFF_save_fm DFF_W4773(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T109));
DFF_save_fm DFF_W4774(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T119));
DFF_save_fm DFF_W4775(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T129));
DFF_save_fm DFF_W4776(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T209));
DFF_save_fm DFF_W4777(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T219));
DFF_save_fm DFF_W4778(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T229));
DFF_save_fm DFF_W4779(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T00A));
DFF_save_fm DFF_W4780(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T01A));
DFF_save_fm DFF_W4781(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T02A));
DFF_save_fm DFF_W4782(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T10A));
DFF_save_fm DFF_W4783(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T11A));
DFF_save_fm DFF_W4784(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T12A));
DFF_save_fm DFF_W4785(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T20A));
DFF_save_fm DFF_W4786(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T21A));
DFF_save_fm DFF_W4787(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T22A));
DFF_save_fm DFF_W4788(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T00B));
DFF_save_fm DFF_W4789(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T01B));
DFF_save_fm DFF_W4790(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T02B));
DFF_save_fm DFF_W4791(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T10B));
DFF_save_fm DFF_W4792(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T11B));
DFF_save_fm DFF_W4793(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T12B));
DFF_save_fm DFF_W4794(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T20B));
DFF_save_fm DFF_W4795(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T21B));
DFF_save_fm DFF_W4796(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T22B));
DFF_save_fm DFF_W4797(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T00C));
DFF_save_fm DFF_W4798(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T01C));
DFF_save_fm DFF_W4799(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T02C));
DFF_save_fm DFF_W4800(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T10C));
DFF_save_fm DFF_W4801(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T11C));
DFF_save_fm DFF_W4802(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T12C));
DFF_save_fm DFF_W4803(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T20C));
DFF_save_fm DFF_W4804(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T21C));
DFF_save_fm DFF_W4805(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T22C));
DFF_save_fm DFF_W4806(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T00D));
DFF_save_fm DFF_W4807(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T01D));
DFF_save_fm DFF_W4808(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T02D));
DFF_save_fm DFF_W4809(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T10D));
DFF_save_fm DFF_W4810(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T11D));
DFF_save_fm DFF_W4811(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T12D));
DFF_save_fm DFF_W4812(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T20D));
DFF_save_fm DFF_W4813(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T21D));
DFF_save_fm DFF_W4814(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T22D));
DFF_save_fm DFF_W4815(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T00E));
DFF_save_fm DFF_W4816(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T01E));
DFF_save_fm DFF_W4817(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T02E));
DFF_save_fm DFF_W4818(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T10E));
DFF_save_fm DFF_W4819(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T11E));
DFF_save_fm DFF_W4820(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T12E));
DFF_save_fm DFF_W4821(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T20E));
DFF_save_fm DFF_W4822(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T21E));
DFF_save_fm DFF_W4823(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T22E));
DFF_save_fm DFF_W4824(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T00F));
DFF_save_fm DFF_W4825(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T01F));
DFF_save_fm DFF_W4826(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T02F));
DFF_save_fm DFF_W4827(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T10F));
DFF_save_fm DFF_W4828(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T11F));
DFF_save_fm DFF_W4829(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T12F));
DFF_save_fm DFF_W4830(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2T20F));
DFF_save_fm DFF_W4831(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T21F));
DFF_save_fm DFF_W4832(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2T22F));
DFF_save_fm DFF_W4833(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U000));
DFF_save_fm DFF_W4834(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U010));
DFF_save_fm DFF_W4835(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U020));
DFF_save_fm DFF_W4836(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U100));
DFF_save_fm DFF_W4837(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U110));
DFF_save_fm DFF_W4838(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U120));
DFF_save_fm DFF_W4839(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U200));
DFF_save_fm DFF_W4840(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U210));
DFF_save_fm DFF_W4841(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U220));
DFF_save_fm DFF_W4842(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U001));
DFF_save_fm DFF_W4843(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U011));
DFF_save_fm DFF_W4844(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U021));
DFF_save_fm DFF_W4845(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U101));
DFF_save_fm DFF_W4846(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U111));
DFF_save_fm DFF_W4847(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U121));
DFF_save_fm DFF_W4848(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U201));
DFF_save_fm DFF_W4849(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U211));
DFF_save_fm DFF_W4850(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U221));
DFF_save_fm DFF_W4851(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U002));
DFF_save_fm DFF_W4852(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U012));
DFF_save_fm DFF_W4853(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U022));
DFF_save_fm DFF_W4854(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U102));
DFF_save_fm DFF_W4855(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U112));
DFF_save_fm DFF_W4856(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U122));
DFF_save_fm DFF_W4857(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U202));
DFF_save_fm DFF_W4858(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U212));
DFF_save_fm DFF_W4859(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U222));
DFF_save_fm DFF_W4860(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U003));
DFF_save_fm DFF_W4861(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U013));
DFF_save_fm DFF_W4862(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U023));
DFF_save_fm DFF_W4863(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U103));
DFF_save_fm DFF_W4864(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U113));
DFF_save_fm DFF_W4865(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U123));
DFF_save_fm DFF_W4866(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U203));
DFF_save_fm DFF_W4867(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U213));
DFF_save_fm DFF_W4868(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U223));
DFF_save_fm DFF_W4869(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U004));
DFF_save_fm DFF_W4870(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U014));
DFF_save_fm DFF_W4871(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U024));
DFF_save_fm DFF_W4872(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U104));
DFF_save_fm DFF_W4873(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U114));
DFF_save_fm DFF_W4874(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U124));
DFF_save_fm DFF_W4875(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U204));
DFF_save_fm DFF_W4876(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U214));
DFF_save_fm DFF_W4877(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U224));
DFF_save_fm DFF_W4878(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U005));
DFF_save_fm DFF_W4879(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U015));
DFF_save_fm DFF_W4880(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U025));
DFF_save_fm DFF_W4881(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U105));
DFF_save_fm DFF_W4882(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U115));
DFF_save_fm DFF_W4883(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U125));
DFF_save_fm DFF_W4884(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U205));
DFF_save_fm DFF_W4885(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U215));
DFF_save_fm DFF_W4886(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U225));
DFF_save_fm DFF_W4887(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U006));
DFF_save_fm DFF_W4888(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U016));
DFF_save_fm DFF_W4889(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U026));
DFF_save_fm DFF_W4890(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U106));
DFF_save_fm DFF_W4891(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U116));
DFF_save_fm DFF_W4892(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U126));
DFF_save_fm DFF_W4893(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U206));
DFF_save_fm DFF_W4894(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U216));
DFF_save_fm DFF_W4895(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U226));
DFF_save_fm DFF_W4896(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U007));
DFF_save_fm DFF_W4897(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U017));
DFF_save_fm DFF_W4898(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U027));
DFF_save_fm DFF_W4899(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U107));
DFF_save_fm DFF_W4900(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U117));
DFF_save_fm DFF_W4901(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U127));
DFF_save_fm DFF_W4902(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U207));
DFF_save_fm DFF_W4903(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U217));
DFF_save_fm DFF_W4904(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U227));
DFF_save_fm DFF_W4905(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U008));
DFF_save_fm DFF_W4906(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U018));
DFF_save_fm DFF_W4907(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U028));
DFF_save_fm DFF_W4908(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U108));
DFF_save_fm DFF_W4909(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U118));
DFF_save_fm DFF_W4910(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U128));
DFF_save_fm DFF_W4911(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U208));
DFF_save_fm DFF_W4912(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U218));
DFF_save_fm DFF_W4913(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U228));
DFF_save_fm DFF_W4914(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U009));
DFF_save_fm DFF_W4915(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U019));
DFF_save_fm DFF_W4916(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U029));
DFF_save_fm DFF_W4917(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U109));
DFF_save_fm DFF_W4918(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U119));
DFF_save_fm DFF_W4919(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U129));
DFF_save_fm DFF_W4920(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U209));
DFF_save_fm DFF_W4921(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U219));
DFF_save_fm DFF_W4922(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U229));
DFF_save_fm DFF_W4923(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U00A));
DFF_save_fm DFF_W4924(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U01A));
DFF_save_fm DFF_W4925(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U02A));
DFF_save_fm DFF_W4926(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U10A));
DFF_save_fm DFF_W4927(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U11A));
DFF_save_fm DFF_W4928(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U12A));
DFF_save_fm DFF_W4929(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U20A));
DFF_save_fm DFF_W4930(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U21A));
DFF_save_fm DFF_W4931(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U22A));
DFF_save_fm DFF_W4932(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U00B));
DFF_save_fm DFF_W4933(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U01B));
DFF_save_fm DFF_W4934(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U02B));
DFF_save_fm DFF_W4935(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U10B));
DFF_save_fm DFF_W4936(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U11B));
DFF_save_fm DFF_W4937(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U12B));
DFF_save_fm DFF_W4938(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U20B));
DFF_save_fm DFF_W4939(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U21B));
DFF_save_fm DFF_W4940(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U22B));
DFF_save_fm DFF_W4941(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U00C));
DFF_save_fm DFF_W4942(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U01C));
DFF_save_fm DFF_W4943(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U02C));
DFF_save_fm DFF_W4944(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U10C));
DFF_save_fm DFF_W4945(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U11C));
DFF_save_fm DFF_W4946(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U12C));
DFF_save_fm DFF_W4947(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U20C));
DFF_save_fm DFF_W4948(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U21C));
DFF_save_fm DFF_W4949(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U22C));
DFF_save_fm DFF_W4950(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U00D));
DFF_save_fm DFF_W4951(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U01D));
DFF_save_fm DFF_W4952(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U02D));
DFF_save_fm DFF_W4953(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U10D));
DFF_save_fm DFF_W4954(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U11D));
DFF_save_fm DFF_W4955(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U12D));
DFF_save_fm DFF_W4956(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U20D));
DFF_save_fm DFF_W4957(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U21D));
DFF_save_fm DFF_W4958(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U22D));
DFF_save_fm DFF_W4959(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U00E));
DFF_save_fm DFF_W4960(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U01E));
DFF_save_fm DFF_W4961(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U02E));
DFF_save_fm DFF_W4962(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U10E));
DFF_save_fm DFF_W4963(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U11E));
DFF_save_fm DFF_W4964(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U12E));
DFF_save_fm DFF_W4965(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U20E));
DFF_save_fm DFF_W4966(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U21E));
DFF_save_fm DFF_W4967(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U22E));
DFF_save_fm DFF_W4968(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U00F));
DFF_save_fm DFF_W4969(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U01F));
DFF_save_fm DFF_W4970(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U02F));
DFF_save_fm DFF_W4971(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U10F));
DFF_save_fm DFF_W4972(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2U11F));
DFF_save_fm DFF_W4973(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U12F));
DFF_save_fm DFF_W4974(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U20F));
DFF_save_fm DFF_W4975(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U21F));
DFF_save_fm DFF_W4976(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2U22F));
DFF_save_fm DFF_W4977(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V000));
DFF_save_fm DFF_W4978(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V010));
DFF_save_fm DFF_W4979(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V020));
DFF_save_fm DFF_W4980(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V100));
DFF_save_fm DFF_W4981(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V110));
DFF_save_fm DFF_W4982(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V120));
DFF_save_fm DFF_W4983(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V200));
DFF_save_fm DFF_W4984(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V210));
DFF_save_fm DFF_W4985(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V220));
DFF_save_fm DFF_W4986(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V001));
DFF_save_fm DFF_W4987(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V011));
DFF_save_fm DFF_W4988(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V021));
DFF_save_fm DFF_W4989(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V101));
DFF_save_fm DFF_W4990(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V111));
DFF_save_fm DFF_W4991(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V121));
DFF_save_fm DFF_W4992(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V201));
DFF_save_fm DFF_W4993(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V211));
DFF_save_fm DFF_W4994(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V221));
DFF_save_fm DFF_W4995(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V002));
DFF_save_fm DFF_W4996(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V012));
DFF_save_fm DFF_W4997(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V022));
DFF_save_fm DFF_W4998(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V102));
DFF_save_fm DFF_W4999(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V112));
DFF_save_fm DFF_W5000(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V122));
DFF_save_fm DFF_W5001(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V202));
DFF_save_fm DFF_W5002(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V212));
DFF_save_fm DFF_W5003(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V222));
DFF_save_fm DFF_W5004(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V003));
DFF_save_fm DFF_W5005(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V013));
DFF_save_fm DFF_W5006(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V023));
DFF_save_fm DFF_W5007(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V103));
DFF_save_fm DFF_W5008(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V113));
DFF_save_fm DFF_W5009(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V123));
DFF_save_fm DFF_W5010(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V203));
DFF_save_fm DFF_W5011(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V213));
DFF_save_fm DFF_W5012(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V223));
DFF_save_fm DFF_W5013(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V004));
DFF_save_fm DFF_W5014(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V014));
DFF_save_fm DFF_W5015(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V024));
DFF_save_fm DFF_W5016(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V104));
DFF_save_fm DFF_W5017(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V114));
DFF_save_fm DFF_W5018(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V124));
DFF_save_fm DFF_W5019(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V204));
DFF_save_fm DFF_W5020(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V214));
DFF_save_fm DFF_W5021(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V224));
DFF_save_fm DFF_W5022(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V005));
DFF_save_fm DFF_W5023(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V015));
DFF_save_fm DFF_W5024(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V025));
DFF_save_fm DFF_W5025(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V105));
DFF_save_fm DFF_W5026(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V115));
DFF_save_fm DFF_W5027(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V125));
DFF_save_fm DFF_W5028(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V205));
DFF_save_fm DFF_W5029(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V215));
DFF_save_fm DFF_W5030(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V225));
DFF_save_fm DFF_W5031(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V006));
DFF_save_fm DFF_W5032(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V016));
DFF_save_fm DFF_W5033(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V026));
DFF_save_fm DFF_W5034(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V106));
DFF_save_fm DFF_W5035(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V116));
DFF_save_fm DFF_W5036(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V126));
DFF_save_fm DFF_W5037(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V206));
DFF_save_fm DFF_W5038(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V216));
DFF_save_fm DFF_W5039(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V226));
DFF_save_fm DFF_W5040(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V007));
DFF_save_fm DFF_W5041(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V017));
DFF_save_fm DFF_W5042(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V027));
DFF_save_fm DFF_W5043(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V107));
DFF_save_fm DFF_W5044(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V117));
DFF_save_fm DFF_W5045(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V127));
DFF_save_fm DFF_W5046(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V207));
DFF_save_fm DFF_W5047(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V217));
DFF_save_fm DFF_W5048(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V227));
DFF_save_fm DFF_W5049(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V008));
DFF_save_fm DFF_W5050(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V018));
DFF_save_fm DFF_W5051(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V028));
DFF_save_fm DFF_W5052(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V108));
DFF_save_fm DFF_W5053(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V118));
DFF_save_fm DFF_W5054(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V128));
DFF_save_fm DFF_W5055(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V208));
DFF_save_fm DFF_W5056(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V218));
DFF_save_fm DFF_W5057(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V228));
DFF_save_fm DFF_W5058(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V009));
DFF_save_fm DFF_W5059(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V019));
DFF_save_fm DFF_W5060(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V029));
DFF_save_fm DFF_W5061(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V109));
DFF_save_fm DFF_W5062(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V119));
DFF_save_fm DFF_W5063(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V129));
DFF_save_fm DFF_W5064(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V209));
DFF_save_fm DFF_W5065(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V219));
DFF_save_fm DFF_W5066(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V229));
DFF_save_fm DFF_W5067(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V00A));
DFF_save_fm DFF_W5068(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V01A));
DFF_save_fm DFF_W5069(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V02A));
DFF_save_fm DFF_W5070(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V10A));
DFF_save_fm DFF_W5071(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V11A));
DFF_save_fm DFF_W5072(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V12A));
DFF_save_fm DFF_W5073(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V20A));
DFF_save_fm DFF_W5074(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V21A));
DFF_save_fm DFF_W5075(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V22A));
DFF_save_fm DFF_W5076(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V00B));
DFF_save_fm DFF_W5077(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V01B));
DFF_save_fm DFF_W5078(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V02B));
DFF_save_fm DFF_W5079(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V10B));
DFF_save_fm DFF_W5080(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V11B));
DFF_save_fm DFF_W5081(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V12B));
DFF_save_fm DFF_W5082(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V20B));
DFF_save_fm DFF_W5083(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V21B));
DFF_save_fm DFF_W5084(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V22B));
DFF_save_fm DFF_W5085(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V00C));
DFF_save_fm DFF_W5086(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V01C));
DFF_save_fm DFF_W5087(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V02C));
DFF_save_fm DFF_W5088(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V10C));
DFF_save_fm DFF_W5089(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V11C));
DFF_save_fm DFF_W5090(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V12C));
DFF_save_fm DFF_W5091(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V20C));
DFF_save_fm DFF_W5092(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V21C));
DFF_save_fm DFF_W5093(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V22C));
DFF_save_fm DFF_W5094(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V00D));
DFF_save_fm DFF_W5095(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V01D));
DFF_save_fm DFF_W5096(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V02D));
DFF_save_fm DFF_W5097(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V10D));
DFF_save_fm DFF_W5098(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V11D));
DFF_save_fm DFF_W5099(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V12D));
DFF_save_fm DFF_W5100(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V20D));
DFF_save_fm DFF_W5101(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V21D));
DFF_save_fm DFF_W5102(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V22D));
DFF_save_fm DFF_W5103(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V00E));
DFF_save_fm DFF_W5104(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V01E));
DFF_save_fm DFF_W5105(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V02E));
DFF_save_fm DFF_W5106(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V10E));
DFF_save_fm DFF_W5107(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V11E));
DFF_save_fm DFF_W5108(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V12E));
DFF_save_fm DFF_W5109(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V20E));
DFF_save_fm DFF_W5110(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V21E));
DFF_save_fm DFF_W5111(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V22E));
DFF_save_fm DFF_W5112(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V00F));
DFF_save_fm DFF_W5113(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V01F));
DFF_save_fm DFF_W5114(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V02F));
DFF_save_fm DFF_W5115(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V10F));
DFF_save_fm DFF_W5116(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V11F));
DFF_save_fm DFF_W5117(.clk(clk),.rstn(rstn),.reset_value(1),.q(W2V12F));
DFF_save_fm DFF_W5118(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V20F));
DFF_save_fm DFF_W5119(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V21F));
DFF_save_fm DFF_W5120(.clk(clk),.rstn(rstn),.reset_value(0),.q(W2V22F));
ninexnine_unit ninexnine_unit_2964(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20000)
);

ninexnine_unit ninexnine_unit_2965(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21000)
);

ninexnine_unit ninexnine_unit_2966(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22000)
);

ninexnine_unit ninexnine_unit_2967(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23000)
);

ninexnine_unit ninexnine_unit_2968(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24000)
);

ninexnine_unit ninexnine_unit_2969(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25000)
);

ninexnine_unit ninexnine_unit_2970(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26000)
);

ninexnine_unit ninexnine_unit_2971(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27000)
);

ninexnine_unit ninexnine_unit_2972(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W20008),
				.b1(W20018),
				.b2(W20028),
				.b3(W20108),
				.b4(W20118),
				.b5(W20128),
				.b6(W20208),
				.b7(W20218),
				.b8(W20228),
				.c(c28000)
);

ninexnine_unit ninexnine_unit_2973(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W20009),
				.b1(W20019),
				.b2(W20029),
				.b3(W20109),
				.b4(W20119),
				.b5(W20129),
				.b6(W20209),
				.b7(W20219),
				.b8(W20229),
				.c(c29000)
);

ninexnine_unit ninexnine_unit_2974(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2000A),
				.b1(W2001A),
				.b2(W2002A),
				.b3(W2010A),
				.b4(W2011A),
				.b5(W2012A),
				.b6(W2020A),
				.b7(W2021A),
				.b8(W2022A),
				.c(c2A000)
);

ninexnine_unit ninexnine_unit_2975(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2000B),
				.b1(W2001B),
				.b2(W2002B),
				.b3(W2010B),
				.b4(W2011B),
				.b5(W2012B),
				.b6(W2020B),
				.b7(W2021B),
				.b8(W2022B),
				.c(c2B000)
);

ninexnine_unit ninexnine_unit_2976(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2000C),
				.b1(W2001C),
				.b2(W2002C),
				.b3(W2010C),
				.b4(W2011C),
				.b5(W2012C),
				.b6(W2020C),
				.b7(W2021C),
				.b8(W2022C),
				.c(c2C000)
);

ninexnine_unit ninexnine_unit_2977(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2000D),
				.b1(W2001D),
				.b2(W2002D),
				.b3(W2010D),
				.b4(W2011D),
				.b5(W2012D),
				.b6(W2020D),
				.b7(W2021D),
				.b8(W2022D),
				.c(c2D000)
);

ninexnine_unit ninexnine_unit_2978(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2000E),
				.b1(W2001E),
				.b2(W2002E),
				.b3(W2010E),
				.b4(W2011E),
				.b5(W2012E),
				.b6(W2020E),
				.b7(W2021E),
				.b8(W2022E),
				.c(c2E000)
);

ninexnine_unit ninexnine_unit_2979(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2000F),
				.b1(W2001F),
				.b2(W2002F),
				.b3(W2010F),
				.b4(W2011F),
				.b5(W2012F),
				.b6(W2020F),
				.b7(W2021F),
				.b8(W2022F),
				.c(c2F000)
);

assign C2000=c20000+c21000+c22000+c23000+c24000+c25000+c26000+c27000+c28000+c29000+c2A000+c2B000+c2C000+c2D000+c2E000+c2F000;
assign A2000=(C2000>=0)?1:0;

assign P3000=A2000;

ninexnine_unit ninexnine_unit_2980(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20010)
);

ninexnine_unit ninexnine_unit_2981(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21010)
);

ninexnine_unit ninexnine_unit_2982(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22010)
);

ninexnine_unit ninexnine_unit_2983(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23010)
);

ninexnine_unit ninexnine_unit_2984(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24010)
);

ninexnine_unit ninexnine_unit_2985(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25010)
);

ninexnine_unit ninexnine_unit_2986(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26010)
);

ninexnine_unit ninexnine_unit_2987(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27010)
);

ninexnine_unit ninexnine_unit_2988(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W20008),
				.b1(W20018),
				.b2(W20028),
				.b3(W20108),
				.b4(W20118),
				.b5(W20128),
				.b6(W20208),
				.b7(W20218),
				.b8(W20228),
				.c(c28010)
);

ninexnine_unit ninexnine_unit_2989(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W20009),
				.b1(W20019),
				.b2(W20029),
				.b3(W20109),
				.b4(W20119),
				.b5(W20129),
				.b6(W20209),
				.b7(W20219),
				.b8(W20229),
				.c(c29010)
);

ninexnine_unit ninexnine_unit_2990(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2000A),
				.b1(W2001A),
				.b2(W2002A),
				.b3(W2010A),
				.b4(W2011A),
				.b5(W2012A),
				.b6(W2020A),
				.b7(W2021A),
				.b8(W2022A),
				.c(c2A010)
);

ninexnine_unit ninexnine_unit_2991(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2000B),
				.b1(W2001B),
				.b2(W2002B),
				.b3(W2010B),
				.b4(W2011B),
				.b5(W2012B),
				.b6(W2020B),
				.b7(W2021B),
				.b8(W2022B),
				.c(c2B010)
);

ninexnine_unit ninexnine_unit_2992(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2000C),
				.b1(W2001C),
				.b2(W2002C),
				.b3(W2010C),
				.b4(W2011C),
				.b5(W2012C),
				.b6(W2020C),
				.b7(W2021C),
				.b8(W2022C),
				.c(c2C010)
);

ninexnine_unit ninexnine_unit_2993(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2000D),
				.b1(W2001D),
				.b2(W2002D),
				.b3(W2010D),
				.b4(W2011D),
				.b5(W2012D),
				.b6(W2020D),
				.b7(W2021D),
				.b8(W2022D),
				.c(c2D010)
);

ninexnine_unit ninexnine_unit_2994(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2000E),
				.b1(W2001E),
				.b2(W2002E),
				.b3(W2010E),
				.b4(W2011E),
				.b5(W2012E),
				.b6(W2020E),
				.b7(W2021E),
				.b8(W2022E),
				.c(c2E010)
);

ninexnine_unit ninexnine_unit_2995(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2000F),
				.b1(W2001F),
				.b2(W2002F),
				.b3(W2010F),
				.b4(W2011F),
				.b5(W2012F),
				.b6(W2020F),
				.b7(W2021F),
				.b8(W2022F),
				.c(c2F010)
);

assign C2010=c20010+c21010+c22010+c23010+c24010+c25010+c26010+c27010+c28010+c29010+c2A010+c2B010+c2C010+c2D010+c2E010+c2F010;
assign A2010=(C2010>=0)?1:0;

assign P3010=A2010;

ninexnine_unit ninexnine_unit_2996(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20020)
);

ninexnine_unit ninexnine_unit_2997(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21020)
);

ninexnine_unit ninexnine_unit_2998(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22020)
);

ninexnine_unit ninexnine_unit_2999(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23020)
);

ninexnine_unit ninexnine_unit_3000(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24020)
);

ninexnine_unit ninexnine_unit_3001(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25020)
);

ninexnine_unit ninexnine_unit_3002(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26020)
);

ninexnine_unit ninexnine_unit_3003(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27020)
);

ninexnine_unit ninexnine_unit_3004(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W20008),
				.b1(W20018),
				.b2(W20028),
				.b3(W20108),
				.b4(W20118),
				.b5(W20128),
				.b6(W20208),
				.b7(W20218),
				.b8(W20228),
				.c(c28020)
);

ninexnine_unit ninexnine_unit_3005(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W20009),
				.b1(W20019),
				.b2(W20029),
				.b3(W20109),
				.b4(W20119),
				.b5(W20129),
				.b6(W20209),
				.b7(W20219),
				.b8(W20229),
				.c(c29020)
);

ninexnine_unit ninexnine_unit_3006(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2000A),
				.b1(W2001A),
				.b2(W2002A),
				.b3(W2010A),
				.b4(W2011A),
				.b5(W2012A),
				.b6(W2020A),
				.b7(W2021A),
				.b8(W2022A),
				.c(c2A020)
);

ninexnine_unit ninexnine_unit_3007(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2000B),
				.b1(W2001B),
				.b2(W2002B),
				.b3(W2010B),
				.b4(W2011B),
				.b5(W2012B),
				.b6(W2020B),
				.b7(W2021B),
				.b8(W2022B),
				.c(c2B020)
);

ninexnine_unit ninexnine_unit_3008(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2000C),
				.b1(W2001C),
				.b2(W2002C),
				.b3(W2010C),
				.b4(W2011C),
				.b5(W2012C),
				.b6(W2020C),
				.b7(W2021C),
				.b8(W2022C),
				.c(c2C020)
);

ninexnine_unit ninexnine_unit_3009(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2000D),
				.b1(W2001D),
				.b2(W2002D),
				.b3(W2010D),
				.b4(W2011D),
				.b5(W2012D),
				.b6(W2020D),
				.b7(W2021D),
				.b8(W2022D),
				.c(c2D020)
);

ninexnine_unit ninexnine_unit_3010(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2000E),
				.b1(W2001E),
				.b2(W2002E),
				.b3(W2010E),
				.b4(W2011E),
				.b5(W2012E),
				.b6(W2020E),
				.b7(W2021E),
				.b8(W2022E),
				.c(c2E020)
);

ninexnine_unit ninexnine_unit_3011(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2000F),
				.b1(W2001F),
				.b2(W2002F),
				.b3(W2010F),
				.b4(W2011F),
				.b5(W2012F),
				.b6(W2020F),
				.b7(W2021F),
				.b8(W2022F),
				.c(c2F020)
);

assign C2020=c20020+c21020+c22020+c23020+c24020+c25020+c26020+c27020+c28020+c29020+c2A020+c2B020+c2C020+c2D020+c2E020+c2F020;
assign A2020=(C2020>=0)?1:0;

assign P3020=A2020;

ninexnine_unit ninexnine_unit_3012(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20100)
);

ninexnine_unit ninexnine_unit_3013(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21100)
);

ninexnine_unit ninexnine_unit_3014(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22100)
);

ninexnine_unit ninexnine_unit_3015(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23100)
);

ninexnine_unit ninexnine_unit_3016(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24100)
);

ninexnine_unit ninexnine_unit_3017(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25100)
);

ninexnine_unit ninexnine_unit_3018(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26100)
);

ninexnine_unit ninexnine_unit_3019(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27100)
);

ninexnine_unit ninexnine_unit_3020(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W20008),
				.b1(W20018),
				.b2(W20028),
				.b3(W20108),
				.b4(W20118),
				.b5(W20128),
				.b6(W20208),
				.b7(W20218),
				.b8(W20228),
				.c(c28100)
);

ninexnine_unit ninexnine_unit_3021(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W20009),
				.b1(W20019),
				.b2(W20029),
				.b3(W20109),
				.b4(W20119),
				.b5(W20129),
				.b6(W20209),
				.b7(W20219),
				.b8(W20229),
				.c(c29100)
);

ninexnine_unit ninexnine_unit_3022(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2000A),
				.b1(W2001A),
				.b2(W2002A),
				.b3(W2010A),
				.b4(W2011A),
				.b5(W2012A),
				.b6(W2020A),
				.b7(W2021A),
				.b8(W2022A),
				.c(c2A100)
);

ninexnine_unit ninexnine_unit_3023(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2000B),
				.b1(W2001B),
				.b2(W2002B),
				.b3(W2010B),
				.b4(W2011B),
				.b5(W2012B),
				.b6(W2020B),
				.b7(W2021B),
				.b8(W2022B),
				.c(c2B100)
);

ninexnine_unit ninexnine_unit_3024(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2000C),
				.b1(W2001C),
				.b2(W2002C),
				.b3(W2010C),
				.b4(W2011C),
				.b5(W2012C),
				.b6(W2020C),
				.b7(W2021C),
				.b8(W2022C),
				.c(c2C100)
);

ninexnine_unit ninexnine_unit_3025(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2000D),
				.b1(W2001D),
				.b2(W2002D),
				.b3(W2010D),
				.b4(W2011D),
				.b5(W2012D),
				.b6(W2020D),
				.b7(W2021D),
				.b8(W2022D),
				.c(c2D100)
);

ninexnine_unit ninexnine_unit_3026(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2000E),
				.b1(W2001E),
				.b2(W2002E),
				.b3(W2010E),
				.b4(W2011E),
				.b5(W2012E),
				.b6(W2020E),
				.b7(W2021E),
				.b8(W2022E),
				.c(c2E100)
);

ninexnine_unit ninexnine_unit_3027(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2000F),
				.b1(W2001F),
				.b2(W2002F),
				.b3(W2010F),
				.b4(W2011F),
				.b5(W2012F),
				.b6(W2020F),
				.b7(W2021F),
				.b8(W2022F),
				.c(c2F100)
);

assign C2100=c20100+c21100+c22100+c23100+c24100+c25100+c26100+c27100+c28100+c29100+c2A100+c2B100+c2C100+c2D100+c2E100+c2F100;
assign A2100=(C2100>=0)?1:0;

assign P3100=A2100;

ninexnine_unit ninexnine_unit_3028(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20110)
);

ninexnine_unit ninexnine_unit_3029(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21110)
);

ninexnine_unit ninexnine_unit_3030(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22110)
);

ninexnine_unit ninexnine_unit_3031(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23110)
);

ninexnine_unit ninexnine_unit_3032(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24110)
);

ninexnine_unit ninexnine_unit_3033(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25110)
);

ninexnine_unit ninexnine_unit_3034(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26110)
);

ninexnine_unit ninexnine_unit_3035(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27110)
);

ninexnine_unit ninexnine_unit_3036(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W20008),
				.b1(W20018),
				.b2(W20028),
				.b3(W20108),
				.b4(W20118),
				.b5(W20128),
				.b6(W20208),
				.b7(W20218),
				.b8(W20228),
				.c(c28110)
);

ninexnine_unit ninexnine_unit_3037(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W20009),
				.b1(W20019),
				.b2(W20029),
				.b3(W20109),
				.b4(W20119),
				.b5(W20129),
				.b6(W20209),
				.b7(W20219),
				.b8(W20229),
				.c(c29110)
);

ninexnine_unit ninexnine_unit_3038(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2000A),
				.b1(W2001A),
				.b2(W2002A),
				.b3(W2010A),
				.b4(W2011A),
				.b5(W2012A),
				.b6(W2020A),
				.b7(W2021A),
				.b8(W2022A),
				.c(c2A110)
);

ninexnine_unit ninexnine_unit_3039(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2000B),
				.b1(W2001B),
				.b2(W2002B),
				.b3(W2010B),
				.b4(W2011B),
				.b5(W2012B),
				.b6(W2020B),
				.b7(W2021B),
				.b8(W2022B),
				.c(c2B110)
);

ninexnine_unit ninexnine_unit_3040(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2000C),
				.b1(W2001C),
				.b2(W2002C),
				.b3(W2010C),
				.b4(W2011C),
				.b5(W2012C),
				.b6(W2020C),
				.b7(W2021C),
				.b8(W2022C),
				.c(c2C110)
);

ninexnine_unit ninexnine_unit_3041(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2000D),
				.b1(W2001D),
				.b2(W2002D),
				.b3(W2010D),
				.b4(W2011D),
				.b5(W2012D),
				.b6(W2020D),
				.b7(W2021D),
				.b8(W2022D),
				.c(c2D110)
);

ninexnine_unit ninexnine_unit_3042(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2000E),
				.b1(W2001E),
				.b2(W2002E),
				.b3(W2010E),
				.b4(W2011E),
				.b5(W2012E),
				.b6(W2020E),
				.b7(W2021E),
				.b8(W2022E),
				.c(c2E110)
);

ninexnine_unit ninexnine_unit_3043(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2000F),
				.b1(W2001F),
				.b2(W2002F),
				.b3(W2010F),
				.b4(W2011F),
				.b5(W2012F),
				.b6(W2020F),
				.b7(W2021F),
				.b8(W2022F),
				.c(c2F110)
);

assign C2110=c20110+c21110+c22110+c23110+c24110+c25110+c26110+c27110+c28110+c29110+c2A110+c2B110+c2C110+c2D110+c2E110+c2F110;
assign A2110=(C2110>=0)?1:0;

assign P3110=A2110;

ninexnine_unit ninexnine_unit_3044(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20120)
);

ninexnine_unit ninexnine_unit_3045(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21120)
);

ninexnine_unit ninexnine_unit_3046(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22120)
);

ninexnine_unit ninexnine_unit_3047(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23120)
);

ninexnine_unit ninexnine_unit_3048(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24120)
);

ninexnine_unit ninexnine_unit_3049(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25120)
);

ninexnine_unit ninexnine_unit_3050(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26120)
);

ninexnine_unit ninexnine_unit_3051(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27120)
);

ninexnine_unit ninexnine_unit_3052(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W20008),
				.b1(W20018),
				.b2(W20028),
				.b3(W20108),
				.b4(W20118),
				.b5(W20128),
				.b6(W20208),
				.b7(W20218),
				.b8(W20228),
				.c(c28120)
);

ninexnine_unit ninexnine_unit_3053(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W20009),
				.b1(W20019),
				.b2(W20029),
				.b3(W20109),
				.b4(W20119),
				.b5(W20129),
				.b6(W20209),
				.b7(W20219),
				.b8(W20229),
				.c(c29120)
);

ninexnine_unit ninexnine_unit_3054(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2000A),
				.b1(W2001A),
				.b2(W2002A),
				.b3(W2010A),
				.b4(W2011A),
				.b5(W2012A),
				.b6(W2020A),
				.b7(W2021A),
				.b8(W2022A),
				.c(c2A120)
);

ninexnine_unit ninexnine_unit_3055(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2000B),
				.b1(W2001B),
				.b2(W2002B),
				.b3(W2010B),
				.b4(W2011B),
				.b5(W2012B),
				.b6(W2020B),
				.b7(W2021B),
				.b8(W2022B),
				.c(c2B120)
);

ninexnine_unit ninexnine_unit_3056(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2000C),
				.b1(W2001C),
				.b2(W2002C),
				.b3(W2010C),
				.b4(W2011C),
				.b5(W2012C),
				.b6(W2020C),
				.b7(W2021C),
				.b8(W2022C),
				.c(c2C120)
);

ninexnine_unit ninexnine_unit_3057(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2000D),
				.b1(W2001D),
				.b2(W2002D),
				.b3(W2010D),
				.b4(W2011D),
				.b5(W2012D),
				.b6(W2020D),
				.b7(W2021D),
				.b8(W2022D),
				.c(c2D120)
);

ninexnine_unit ninexnine_unit_3058(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2000E),
				.b1(W2001E),
				.b2(W2002E),
				.b3(W2010E),
				.b4(W2011E),
				.b5(W2012E),
				.b6(W2020E),
				.b7(W2021E),
				.b8(W2022E),
				.c(c2E120)
);

ninexnine_unit ninexnine_unit_3059(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2000F),
				.b1(W2001F),
				.b2(W2002F),
				.b3(W2010F),
				.b4(W2011F),
				.b5(W2012F),
				.b6(W2020F),
				.b7(W2021F),
				.b8(W2022F),
				.c(c2F120)
);

assign C2120=c20120+c21120+c22120+c23120+c24120+c25120+c26120+c27120+c28120+c29120+c2A120+c2B120+c2C120+c2D120+c2E120+c2F120;
assign A2120=(C2120>=0)?1:0;

assign P3120=A2120;

ninexnine_unit ninexnine_unit_3060(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20200)
);

ninexnine_unit ninexnine_unit_3061(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21200)
);

ninexnine_unit ninexnine_unit_3062(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22200)
);

ninexnine_unit ninexnine_unit_3063(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23200)
);

ninexnine_unit ninexnine_unit_3064(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24200)
);

ninexnine_unit ninexnine_unit_3065(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25200)
);

ninexnine_unit ninexnine_unit_3066(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26200)
);

ninexnine_unit ninexnine_unit_3067(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27200)
);

ninexnine_unit ninexnine_unit_3068(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W20008),
				.b1(W20018),
				.b2(W20028),
				.b3(W20108),
				.b4(W20118),
				.b5(W20128),
				.b6(W20208),
				.b7(W20218),
				.b8(W20228),
				.c(c28200)
);

ninexnine_unit ninexnine_unit_3069(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W20009),
				.b1(W20019),
				.b2(W20029),
				.b3(W20109),
				.b4(W20119),
				.b5(W20129),
				.b6(W20209),
				.b7(W20219),
				.b8(W20229),
				.c(c29200)
);

ninexnine_unit ninexnine_unit_3070(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2000A),
				.b1(W2001A),
				.b2(W2002A),
				.b3(W2010A),
				.b4(W2011A),
				.b5(W2012A),
				.b6(W2020A),
				.b7(W2021A),
				.b8(W2022A),
				.c(c2A200)
);

ninexnine_unit ninexnine_unit_3071(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2000B),
				.b1(W2001B),
				.b2(W2002B),
				.b3(W2010B),
				.b4(W2011B),
				.b5(W2012B),
				.b6(W2020B),
				.b7(W2021B),
				.b8(W2022B),
				.c(c2B200)
);

ninexnine_unit ninexnine_unit_3072(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2000C),
				.b1(W2001C),
				.b2(W2002C),
				.b3(W2010C),
				.b4(W2011C),
				.b5(W2012C),
				.b6(W2020C),
				.b7(W2021C),
				.b8(W2022C),
				.c(c2C200)
);

ninexnine_unit ninexnine_unit_3073(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2000D),
				.b1(W2001D),
				.b2(W2002D),
				.b3(W2010D),
				.b4(W2011D),
				.b5(W2012D),
				.b6(W2020D),
				.b7(W2021D),
				.b8(W2022D),
				.c(c2D200)
);

ninexnine_unit ninexnine_unit_3074(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2000E),
				.b1(W2001E),
				.b2(W2002E),
				.b3(W2010E),
				.b4(W2011E),
				.b5(W2012E),
				.b6(W2020E),
				.b7(W2021E),
				.b8(W2022E),
				.c(c2E200)
);

ninexnine_unit ninexnine_unit_3075(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2000F),
				.b1(W2001F),
				.b2(W2002F),
				.b3(W2010F),
				.b4(W2011F),
				.b5(W2012F),
				.b6(W2020F),
				.b7(W2021F),
				.b8(W2022F),
				.c(c2F200)
);

assign C2200=c20200+c21200+c22200+c23200+c24200+c25200+c26200+c27200+c28200+c29200+c2A200+c2B200+c2C200+c2D200+c2E200+c2F200;
assign A2200=(C2200>=0)?1:0;

assign P3200=A2200;

ninexnine_unit ninexnine_unit_3076(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20210)
);

ninexnine_unit ninexnine_unit_3077(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21210)
);

ninexnine_unit ninexnine_unit_3078(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22210)
);

ninexnine_unit ninexnine_unit_3079(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23210)
);

ninexnine_unit ninexnine_unit_3080(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24210)
);

ninexnine_unit ninexnine_unit_3081(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25210)
);

ninexnine_unit ninexnine_unit_3082(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26210)
);

ninexnine_unit ninexnine_unit_3083(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27210)
);

ninexnine_unit ninexnine_unit_3084(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W20008),
				.b1(W20018),
				.b2(W20028),
				.b3(W20108),
				.b4(W20118),
				.b5(W20128),
				.b6(W20208),
				.b7(W20218),
				.b8(W20228),
				.c(c28210)
);

ninexnine_unit ninexnine_unit_3085(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W20009),
				.b1(W20019),
				.b2(W20029),
				.b3(W20109),
				.b4(W20119),
				.b5(W20129),
				.b6(W20209),
				.b7(W20219),
				.b8(W20229),
				.c(c29210)
);

ninexnine_unit ninexnine_unit_3086(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2000A),
				.b1(W2001A),
				.b2(W2002A),
				.b3(W2010A),
				.b4(W2011A),
				.b5(W2012A),
				.b6(W2020A),
				.b7(W2021A),
				.b8(W2022A),
				.c(c2A210)
);

ninexnine_unit ninexnine_unit_3087(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2000B),
				.b1(W2001B),
				.b2(W2002B),
				.b3(W2010B),
				.b4(W2011B),
				.b5(W2012B),
				.b6(W2020B),
				.b7(W2021B),
				.b8(W2022B),
				.c(c2B210)
);

ninexnine_unit ninexnine_unit_3088(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2000C),
				.b1(W2001C),
				.b2(W2002C),
				.b3(W2010C),
				.b4(W2011C),
				.b5(W2012C),
				.b6(W2020C),
				.b7(W2021C),
				.b8(W2022C),
				.c(c2C210)
);

ninexnine_unit ninexnine_unit_3089(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2000D),
				.b1(W2001D),
				.b2(W2002D),
				.b3(W2010D),
				.b4(W2011D),
				.b5(W2012D),
				.b6(W2020D),
				.b7(W2021D),
				.b8(W2022D),
				.c(c2D210)
);

ninexnine_unit ninexnine_unit_3090(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2000E),
				.b1(W2001E),
				.b2(W2002E),
				.b3(W2010E),
				.b4(W2011E),
				.b5(W2012E),
				.b6(W2020E),
				.b7(W2021E),
				.b8(W2022E),
				.c(c2E210)
);

ninexnine_unit ninexnine_unit_3091(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2000F),
				.b1(W2001F),
				.b2(W2002F),
				.b3(W2010F),
				.b4(W2011F),
				.b5(W2012F),
				.b6(W2020F),
				.b7(W2021F),
				.b8(W2022F),
				.c(c2F210)
);

assign C2210=c20210+c21210+c22210+c23210+c24210+c25210+c26210+c27210+c28210+c29210+c2A210+c2B210+c2C210+c2D210+c2E210+c2F210;
assign A2210=(C2210>=0)?1:0;

assign P3210=A2210;

ninexnine_unit ninexnine_unit_3092(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W20000),
				.b1(W20010),
				.b2(W20020),
				.b3(W20100),
				.b4(W20110),
				.b5(W20120),
				.b6(W20200),
				.b7(W20210),
				.b8(W20220),
				.c(c20220)
);

ninexnine_unit ninexnine_unit_3093(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W20001),
				.b1(W20011),
				.b2(W20021),
				.b3(W20101),
				.b4(W20111),
				.b5(W20121),
				.b6(W20201),
				.b7(W20211),
				.b8(W20221),
				.c(c21220)
);

ninexnine_unit ninexnine_unit_3094(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W20002),
				.b1(W20012),
				.b2(W20022),
				.b3(W20102),
				.b4(W20112),
				.b5(W20122),
				.b6(W20202),
				.b7(W20212),
				.b8(W20222),
				.c(c22220)
);

ninexnine_unit ninexnine_unit_3095(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W20003),
				.b1(W20013),
				.b2(W20023),
				.b3(W20103),
				.b4(W20113),
				.b5(W20123),
				.b6(W20203),
				.b7(W20213),
				.b8(W20223),
				.c(c23220)
);

ninexnine_unit ninexnine_unit_3096(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W20004),
				.b1(W20014),
				.b2(W20024),
				.b3(W20104),
				.b4(W20114),
				.b5(W20124),
				.b6(W20204),
				.b7(W20214),
				.b8(W20224),
				.c(c24220)
);

ninexnine_unit ninexnine_unit_3097(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W20005),
				.b1(W20015),
				.b2(W20025),
				.b3(W20105),
				.b4(W20115),
				.b5(W20125),
				.b6(W20205),
				.b7(W20215),
				.b8(W20225),
				.c(c25220)
);

ninexnine_unit ninexnine_unit_3098(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W20006),
				.b1(W20016),
				.b2(W20026),
				.b3(W20106),
				.b4(W20116),
				.b5(W20126),
				.b6(W20206),
				.b7(W20216),
				.b8(W20226),
				.c(c26220)
);

ninexnine_unit ninexnine_unit_3099(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W20007),
				.b1(W20017),
				.b2(W20027),
				.b3(W20107),
				.b4(W20117),
				.b5(W20127),
				.b6(W20207),
				.b7(W20217),
				.b8(W20227),
				.c(c27220)
);

ninexnine_unit ninexnine_unit_3100(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W20008),
				.b1(W20018),
				.b2(W20028),
				.b3(W20108),
				.b4(W20118),
				.b5(W20128),
				.b6(W20208),
				.b7(W20218),
				.b8(W20228),
				.c(c28220)
);

ninexnine_unit ninexnine_unit_3101(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W20009),
				.b1(W20019),
				.b2(W20029),
				.b3(W20109),
				.b4(W20119),
				.b5(W20129),
				.b6(W20209),
				.b7(W20219),
				.b8(W20229),
				.c(c29220)
);

ninexnine_unit ninexnine_unit_3102(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2000A),
				.b1(W2001A),
				.b2(W2002A),
				.b3(W2010A),
				.b4(W2011A),
				.b5(W2012A),
				.b6(W2020A),
				.b7(W2021A),
				.b8(W2022A),
				.c(c2A220)
);

ninexnine_unit ninexnine_unit_3103(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2000B),
				.b1(W2001B),
				.b2(W2002B),
				.b3(W2010B),
				.b4(W2011B),
				.b5(W2012B),
				.b6(W2020B),
				.b7(W2021B),
				.b8(W2022B),
				.c(c2B220)
);

ninexnine_unit ninexnine_unit_3104(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2000C),
				.b1(W2001C),
				.b2(W2002C),
				.b3(W2010C),
				.b4(W2011C),
				.b5(W2012C),
				.b6(W2020C),
				.b7(W2021C),
				.b8(W2022C),
				.c(c2C220)
);

ninexnine_unit ninexnine_unit_3105(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2000D),
				.b1(W2001D),
				.b2(W2002D),
				.b3(W2010D),
				.b4(W2011D),
				.b5(W2012D),
				.b6(W2020D),
				.b7(W2021D),
				.b8(W2022D),
				.c(c2D220)
);

ninexnine_unit ninexnine_unit_3106(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2000E),
				.b1(W2001E),
				.b2(W2002E),
				.b3(W2010E),
				.b4(W2011E),
				.b5(W2012E),
				.b6(W2020E),
				.b7(W2021E),
				.b8(W2022E),
				.c(c2E220)
);

ninexnine_unit ninexnine_unit_3107(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2000F),
				.b1(W2001F),
				.b2(W2002F),
				.b3(W2010F),
				.b4(W2011F),
				.b5(W2012F),
				.b6(W2020F),
				.b7(W2021F),
				.b8(W2022F),
				.c(c2F220)
);

assign C2220=c20220+c21220+c22220+c23220+c24220+c25220+c26220+c27220+c28220+c29220+c2A220+c2B220+c2C220+c2D220+c2E220+c2F220;
assign A2220=(C2220>=0)?1:0;

assign P3220=A2220;

ninexnine_unit ninexnine_unit_3108(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20001)
);

ninexnine_unit ninexnine_unit_3109(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21001)
);

ninexnine_unit ninexnine_unit_3110(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22001)
);

ninexnine_unit ninexnine_unit_3111(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23001)
);

ninexnine_unit ninexnine_unit_3112(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24001)
);

ninexnine_unit ninexnine_unit_3113(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25001)
);

ninexnine_unit ninexnine_unit_3114(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26001)
);

ninexnine_unit ninexnine_unit_3115(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27001)
);

ninexnine_unit ninexnine_unit_3116(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W21008),
				.b1(W21018),
				.b2(W21028),
				.b3(W21108),
				.b4(W21118),
				.b5(W21128),
				.b6(W21208),
				.b7(W21218),
				.b8(W21228),
				.c(c28001)
);

ninexnine_unit ninexnine_unit_3117(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W21009),
				.b1(W21019),
				.b2(W21029),
				.b3(W21109),
				.b4(W21119),
				.b5(W21129),
				.b6(W21209),
				.b7(W21219),
				.b8(W21229),
				.c(c29001)
);

ninexnine_unit ninexnine_unit_3118(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2100A),
				.b1(W2101A),
				.b2(W2102A),
				.b3(W2110A),
				.b4(W2111A),
				.b5(W2112A),
				.b6(W2120A),
				.b7(W2121A),
				.b8(W2122A),
				.c(c2A001)
);

ninexnine_unit ninexnine_unit_3119(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2100B),
				.b1(W2101B),
				.b2(W2102B),
				.b3(W2110B),
				.b4(W2111B),
				.b5(W2112B),
				.b6(W2120B),
				.b7(W2121B),
				.b8(W2122B),
				.c(c2B001)
);

ninexnine_unit ninexnine_unit_3120(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2100C),
				.b1(W2101C),
				.b2(W2102C),
				.b3(W2110C),
				.b4(W2111C),
				.b5(W2112C),
				.b6(W2120C),
				.b7(W2121C),
				.b8(W2122C),
				.c(c2C001)
);

ninexnine_unit ninexnine_unit_3121(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2100D),
				.b1(W2101D),
				.b2(W2102D),
				.b3(W2110D),
				.b4(W2111D),
				.b5(W2112D),
				.b6(W2120D),
				.b7(W2121D),
				.b8(W2122D),
				.c(c2D001)
);

ninexnine_unit ninexnine_unit_3122(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2100E),
				.b1(W2101E),
				.b2(W2102E),
				.b3(W2110E),
				.b4(W2111E),
				.b5(W2112E),
				.b6(W2120E),
				.b7(W2121E),
				.b8(W2122E),
				.c(c2E001)
);

ninexnine_unit ninexnine_unit_3123(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2100F),
				.b1(W2101F),
				.b2(W2102F),
				.b3(W2110F),
				.b4(W2111F),
				.b5(W2112F),
				.b6(W2120F),
				.b7(W2121F),
				.b8(W2122F),
				.c(c2F001)
);

assign C2001=c20001+c21001+c22001+c23001+c24001+c25001+c26001+c27001+c28001+c29001+c2A001+c2B001+c2C001+c2D001+c2E001+c2F001;
assign A2001=(C2001>=0)?1:0;

assign P3001=A2001;

ninexnine_unit ninexnine_unit_3124(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20011)
);

ninexnine_unit ninexnine_unit_3125(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21011)
);

ninexnine_unit ninexnine_unit_3126(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22011)
);

ninexnine_unit ninexnine_unit_3127(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23011)
);

ninexnine_unit ninexnine_unit_3128(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24011)
);

ninexnine_unit ninexnine_unit_3129(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25011)
);

ninexnine_unit ninexnine_unit_3130(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26011)
);

ninexnine_unit ninexnine_unit_3131(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27011)
);

ninexnine_unit ninexnine_unit_3132(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W21008),
				.b1(W21018),
				.b2(W21028),
				.b3(W21108),
				.b4(W21118),
				.b5(W21128),
				.b6(W21208),
				.b7(W21218),
				.b8(W21228),
				.c(c28011)
);

ninexnine_unit ninexnine_unit_3133(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W21009),
				.b1(W21019),
				.b2(W21029),
				.b3(W21109),
				.b4(W21119),
				.b5(W21129),
				.b6(W21209),
				.b7(W21219),
				.b8(W21229),
				.c(c29011)
);

ninexnine_unit ninexnine_unit_3134(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2100A),
				.b1(W2101A),
				.b2(W2102A),
				.b3(W2110A),
				.b4(W2111A),
				.b5(W2112A),
				.b6(W2120A),
				.b7(W2121A),
				.b8(W2122A),
				.c(c2A011)
);

ninexnine_unit ninexnine_unit_3135(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2100B),
				.b1(W2101B),
				.b2(W2102B),
				.b3(W2110B),
				.b4(W2111B),
				.b5(W2112B),
				.b6(W2120B),
				.b7(W2121B),
				.b8(W2122B),
				.c(c2B011)
);

ninexnine_unit ninexnine_unit_3136(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2100C),
				.b1(W2101C),
				.b2(W2102C),
				.b3(W2110C),
				.b4(W2111C),
				.b5(W2112C),
				.b6(W2120C),
				.b7(W2121C),
				.b8(W2122C),
				.c(c2C011)
);

ninexnine_unit ninexnine_unit_3137(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2100D),
				.b1(W2101D),
				.b2(W2102D),
				.b3(W2110D),
				.b4(W2111D),
				.b5(W2112D),
				.b6(W2120D),
				.b7(W2121D),
				.b8(W2122D),
				.c(c2D011)
);

ninexnine_unit ninexnine_unit_3138(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2100E),
				.b1(W2101E),
				.b2(W2102E),
				.b3(W2110E),
				.b4(W2111E),
				.b5(W2112E),
				.b6(W2120E),
				.b7(W2121E),
				.b8(W2122E),
				.c(c2E011)
);

ninexnine_unit ninexnine_unit_3139(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2100F),
				.b1(W2101F),
				.b2(W2102F),
				.b3(W2110F),
				.b4(W2111F),
				.b5(W2112F),
				.b6(W2120F),
				.b7(W2121F),
				.b8(W2122F),
				.c(c2F011)
);

assign C2011=c20011+c21011+c22011+c23011+c24011+c25011+c26011+c27011+c28011+c29011+c2A011+c2B011+c2C011+c2D011+c2E011+c2F011;
assign A2011=(C2011>=0)?1:0;

assign P3011=A2011;

ninexnine_unit ninexnine_unit_3140(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20021)
);

ninexnine_unit ninexnine_unit_3141(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21021)
);

ninexnine_unit ninexnine_unit_3142(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22021)
);

ninexnine_unit ninexnine_unit_3143(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23021)
);

ninexnine_unit ninexnine_unit_3144(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24021)
);

ninexnine_unit ninexnine_unit_3145(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25021)
);

ninexnine_unit ninexnine_unit_3146(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26021)
);

ninexnine_unit ninexnine_unit_3147(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27021)
);

ninexnine_unit ninexnine_unit_3148(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W21008),
				.b1(W21018),
				.b2(W21028),
				.b3(W21108),
				.b4(W21118),
				.b5(W21128),
				.b6(W21208),
				.b7(W21218),
				.b8(W21228),
				.c(c28021)
);

ninexnine_unit ninexnine_unit_3149(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W21009),
				.b1(W21019),
				.b2(W21029),
				.b3(W21109),
				.b4(W21119),
				.b5(W21129),
				.b6(W21209),
				.b7(W21219),
				.b8(W21229),
				.c(c29021)
);

ninexnine_unit ninexnine_unit_3150(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2100A),
				.b1(W2101A),
				.b2(W2102A),
				.b3(W2110A),
				.b4(W2111A),
				.b5(W2112A),
				.b6(W2120A),
				.b7(W2121A),
				.b8(W2122A),
				.c(c2A021)
);

ninexnine_unit ninexnine_unit_3151(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2100B),
				.b1(W2101B),
				.b2(W2102B),
				.b3(W2110B),
				.b4(W2111B),
				.b5(W2112B),
				.b6(W2120B),
				.b7(W2121B),
				.b8(W2122B),
				.c(c2B021)
);

ninexnine_unit ninexnine_unit_3152(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2100C),
				.b1(W2101C),
				.b2(W2102C),
				.b3(W2110C),
				.b4(W2111C),
				.b5(W2112C),
				.b6(W2120C),
				.b7(W2121C),
				.b8(W2122C),
				.c(c2C021)
);

ninexnine_unit ninexnine_unit_3153(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2100D),
				.b1(W2101D),
				.b2(W2102D),
				.b3(W2110D),
				.b4(W2111D),
				.b5(W2112D),
				.b6(W2120D),
				.b7(W2121D),
				.b8(W2122D),
				.c(c2D021)
);

ninexnine_unit ninexnine_unit_3154(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2100E),
				.b1(W2101E),
				.b2(W2102E),
				.b3(W2110E),
				.b4(W2111E),
				.b5(W2112E),
				.b6(W2120E),
				.b7(W2121E),
				.b8(W2122E),
				.c(c2E021)
);

ninexnine_unit ninexnine_unit_3155(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2100F),
				.b1(W2101F),
				.b2(W2102F),
				.b3(W2110F),
				.b4(W2111F),
				.b5(W2112F),
				.b6(W2120F),
				.b7(W2121F),
				.b8(W2122F),
				.c(c2F021)
);

assign C2021=c20021+c21021+c22021+c23021+c24021+c25021+c26021+c27021+c28021+c29021+c2A021+c2B021+c2C021+c2D021+c2E021+c2F021;
assign A2021=(C2021>=0)?1:0;

assign P3021=A2021;

ninexnine_unit ninexnine_unit_3156(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20101)
);

ninexnine_unit ninexnine_unit_3157(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21101)
);

ninexnine_unit ninexnine_unit_3158(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22101)
);

ninexnine_unit ninexnine_unit_3159(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23101)
);

ninexnine_unit ninexnine_unit_3160(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24101)
);

ninexnine_unit ninexnine_unit_3161(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25101)
);

ninexnine_unit ninexnine_unit_3162(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26101)
);

ninexnine_unit ninexnine_unit_3163(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27101)
);

ninexnine_unit ninexnine_unit_3164(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W21008),
				.b1(W21018),
				.b2(W21028),
				.b3(W21108),
				.b4(W21118),
				.b5(W21128),
				.b6(W21208),
				.b7(W21218),
				.b8(W21228),
				.c(c28101)
);

ninexnine_unit ninexnine_unit_3165(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W21009),
				.b1(W21019),
				.b2(W21029),
				.b3(W21109),
				.b4(W21119),
				.b5(W21129),
				.b6(W21209),
				.b7(W21219),
				.b8(W21229),
				.c(c29101)
);

ninexnine_unit ninexnine_unit_3166(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2100A),
				.b1(W2101A),
				.b2(W2102A),
				.b3(W2110A),
				.b4(W2111A),
				.b5(W2112A),
				.b6(W2120A),
				.b7(W2121A),
				.b8(W2122A),
				.c(c2A101)
);

ninexnine_unit ninexnine_unit_3167(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2100B),
				.b1(W2101B),
				.b2(W2102B),
				.b3(W2110B),
				.b4(W2111B),
				.b5(W2112B),
				.b6(W2120B),
				.b7(W2121B),
				.b8(W2122B),
				.c(c2B101)
);

ninexnine_unit ninexnine_unit_3168(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2100C),
				.b1(W2101C),
				.b2(W2102C),
				.b3(W2110C),
				.b4(W2111C),
				.b5(W2112C),
				.b6(W2120C),
				.b7(W2121C),
				.b8(W2122C),
				.c(c2C101)
);

ninexnine_unit ninexnine_unit_3169(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2100D),
				.b1(W2101D),
				.b2(W2102D),
				.b3(W2110D),
				.b4(W2111D),
				.b5(W2112D),
				.b6(W2120D),
				.b7(W2121D),
				.b8(W2122D),
				.c(c2D101)
);

ninexnine_unit ninexnine_unit_3170(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2100E),
				.b1(W2101E),
				.b2(W2102E),
				.b3(W2110E),
				.b4(W2111E),
				.b5(W2112E),
				.b6(W2120E),
				.b7(W2121E),
				.b8(W2122E),
				.c(c2E101)
);

ninexnine_unit ninexnine_unit_3171(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2100F),
				.b1(W2101F),
				.b2(W2102F),
				.b3(W2110F),
				.b4(W2111F),
				.b5(W2112F),
				.b6(W2120F),
				.b7(W2121F),
				.b8(W2122F),
				.c(c2F101)
);

assign C2101=c20101+c21101+c22101+c23101+c24101+c25101+c26101+c27101+c28101+c29101+c2A101+c2B101+c2C101+c2D101+c2E101+c2F101;
assign A2101=(C2101>=0)?1:0;

assign P3101=A2101;

ninexnine_unit ninexnine_unit_3172(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20111)
);

ninexnine_unit ninexnine_unit_3173(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21111)
);

ninexnine_unit ninexnine_unit_3174(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22111)
);

ninexnine_unit ninexnine_unit_3175(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23111)
);

ninexnine_unit ninexnine_unit_3176(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24111)
);

ninexnine_unit ninexnine_unit_3177(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25111)
);

ninexnine_unit ninexnine_unit_3178(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26111)
);

ninexnine_unit ninexnine_unit_3179(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27111)
);

ninexnine_unit ninexnine_unit_3180(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W21008),
				.b1(W21018),
				.b2(W21028),
				.b3(W21108),
				.b4(W21118),
				.b5(W21128),
				.b6(W21208),
				.b7(W21218),
				.b8(W21228),
				.c(c28111)
);

ninexnine_unit ninexnine_unit_3181(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W21009),
				.b1(W21019),
				.b2(W21029),
				.b3(W21109),
				.b4(W21119),
				.b5(W21129),
				.b6(W21209),
				.b7(W21219),
				.b8(W21229),
				.c(c29111)
);

ninexnine_unit ninexnine_unit_3182(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2100A),
				.b1(W2101A),
				.b2(W2102A),
				.b3(W2110A),
				.b4(W2111A),
				.b5(W2112A),
				.b6(W2120A),
				.b7(W2121A),
				.b8(W2122A),
				.c(c2A111)
);

ninexnine_unit ninexnine_unit_3183(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2100B),
				.b1(W2101B),
				.b2(W2102B),
				.b3(W2110B),
				.b4(W2111B),
				.b5(W2112B),
				.b6(W2120B),
				.b7(W2121B),
				.b8(W2122B),
				.c(c2B111)
);

ninexnine_unit ninexnine_unit_3184(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2100C),
				.b1(W2101C),
				.b2(W2102C),
				.b3(W2110C),
				.b4(W2111C),
				.b5(W2112C),
				.b6(W2120C),
				.b7(W2121C),
				.b8(W2122C),
				.c(c2C111)
);

ninexnine_unit ninexnine_unit_3185(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2100D),
				.b1(W2101D),
				.b2(W2102D),
				.b3(W2110D),
				.b4(W2111D),
				.b5(W2112D),
				.b6(W2120D),
				.b7(W2121D),
				.b8(W2122D),
				.c(c2D111)
);

ninexnine_unit ninexnine_unit_3186(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2100E),
				.b1(W2101E),
				.b2(W2102E),
				.b3(W2110E),
				.b4(W2111E),
				.b5(W2112E),
				.b6(W2120E),
				.b7(W2121E),
				.b8(W2122E),
				.c(c2E111)
);

ninexnine_unit ninexnine_unit_3187(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2100F),
				.b1(W2101F),
				.b2(W2102F),
				.b3(W2110F),
				.b4(W2111F),
				.b5(W2112F),
				.b6(W2120F),
				.b7(W2121F),
				.b8(W2122F),
				.c(c2F111)
);

assign C2111=c20111+c21111+c22111+c23111+c24111+c25111+c26111+c27111+c28111+c29111+c2A111+c2B111+c2C111+c2D111+c2E111+c2F111;
assign A2111=(C2111>=0)?1:0;

assign P3111=A2111;

ninexnine_unit ninexnine_unit_3188(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20121)
);

ninexnine_unit ninexnine_unit_3189(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21121)
);

ninexnine_unit ninexnine_unit_3190(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22121)
);

ninexnine_unit ninexnine_unit_3191(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23121)
);

ninexnine_unit ninexnine_unit_3192(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24121)
);

ninexnine_unit ninexnine_unit_3193(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25121)
);

ninexnine_unit ninexnine_unit_3194(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26121)
);

ninexnine_unit ninexnine_unit_3195(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27121)
);

ninexnine_unit ninexnine_unit_3196(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W21008),
				.b1(W21018),
				.b2(W21028),
				.b3(W21108),
				.b4(W21118),
				.b5(W21128),
				.b6(W21208),
				.b7(W21218),
				.b8(W21228),
				.c(c28121)
);

ninexnine_unit ninexnine_unit_3197(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W21009),
				.b1(W21019),
				.b2(W21029),
				.b3(W21109),
				.b4(W21119),
				.b5(W21129),
				.b6(W21209),
				.b7(W21219),
				.b8(W21229),
				.c(c29121)
);

ninexnine_unit ninexnine_unit_3198(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2100A),
				.b1(W2101A),
				.b2(W2102A),
				.b3(W2110A),
				.b4(W2111A),
				.b5(W2112A),
				.b6(W2120A),
				.b7(W2121A),
				.b8(W2122A),
				.c(c2A121)
);

ninexnine_unit ninexnine_unit_3199(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2100B),
				.b1(W2101B),
				.b2(W2102B),
				.b3(W2110B),
				.b4(W2111B),
				.b5(W2112B),
				.b6(W2120B),
				.b7(W2121B),
				.b8(W2122B),
				.c(c2B121)
);

ninexnine_unit ninexnine_unit_3200(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2100C),
				.b1(W2101C),
				.b2(W2102C),
				.b3(W2110C),
				.b4(W2111C),
				.b5(W2112C),
				.b6(W2120C),
				.b7(W2121C),
				.b8(W2122C),
				.c(c2C121)
);

ninexnine_unit ninexnine_unit_3201(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2100D),
				.b1(W2101D),
				.b2(W2102D),
				.b3(W2110D),
				.b4(W2111D),
				.b5(W2112D),
				.b6(W2120D),
				.b7(W2121D),
				.b8(W2122D),
				.c(c2D121)
);

ninexnine_unit ninexnine_unit_3202(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2100E),
				.b1(W2101E),
				.b2(W2102E),
				.b3(W2110E),
				.b4(W2111E),
				.b5(W2112E),
				.b6(W2120E),
				.b7(W2121E),
				.b8(W2122E),
				.c(c2E121)
);

ninexnine_unit ninexnine_unit_3203(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2100F),
				.b1(W2101F),
				.b2(W2102F),
				.b3(W2110F),
				.b4(W2111F),
				.b5(W2112F),
				.b6(W2120F),
				.b7(W2121F),
				.b8(W2122F),
				.c(c2F121)
);

assign C2121=c20121+c21121+c22121+c23121+c24121+c25121+c26121+c27121+c28121+c29121+c2A121+c2B121+c2C121+c2D121+c2E121+c2F121;
assign A2121=(C2121>=0)?1:0;

assign P3121=A2121;

ninexnine_unit ninexnine_unit_3204(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20201)
);

ninexnine_unit ninexnine_unit_3205(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21201)
);

ninexnine_unit ninexnine_unit_3206(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22201)
);

ninexnine_unit ninexnine_unit_3207(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23201)
);

ninexnine_unit ninexnine_unit_3208(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24201)
);

ninexnine_unit ninexnine_unit_3209(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25201)
);

ninexnine_unit ninexnine_unit_3210(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26201)
);

ninexnine_unit ninexnine_unit_3211(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27201)
);

ninexnine_unit ninexnine_unit_3212(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W21008),
				.b1(W21018),
				.b2(W21028),
				.b3(W21108),
				.b4(W21118),
				.b5(W21128),
				.b6(W21208),
				.b7(W21218),
				.b8(W21228),
				.c(c28201)
);

ninexnine_unit ninexnine_unit_3213(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W21009),
				.b1(W21019),
				.b2(W21029),
				.b3(W21109),
				.b4(W21119),
				.b5(W21129),
				.b6(W21209),
				.b7(W21219),
				.b8(W21229),
				.c(c29201)
);

ninexnine_unit ninexnine_unit_3214(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2100A),
				.b1(W2101A),
				.b2(W2102A),
				.b3(W2110A),
				.b4(W2111A),
				.b5(W2112A),
				.b6(W2120A),
				.b7(W2121A),
				.b8(W2122A),
				.c(c2A201)
);

ninexnine_unit ninexnine_unit_3215(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2100B),
				.b1(W2101B),
				.b2(W2102B),
				.b3(W2110B),
				.b4(W2111B),
				.b5(W2112B),
				.b6(W2120B),
				.b7(W2121B),
				.b8(W2122B),
				.c(c2B201)
);

ninexnine_unit ninexnine_unit_3216(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2100C),
				.b1(W2101C),
				.b2(W2102C),
				.b3(W2110C),
				.b4(W2111C),
				.b5(W2112C),
				.b6(W2120C),
				.b7(W2121C),
				.b8(W2122C),
				.c(c2C201)
);

ninexnine_unit ninexnine_unit_3217(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2100D),
				.b1(W2101D),
				.b2(W2102D),
				.b3(W2110D),
				.b4(W2111D),
				.b5(W2112D),
				.b6(W2120D),
				.b7(W2121D),
				.b8(W2122D),
				.c(c2D201)
);

ninexnine_unit ninexnine_unit_3218(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2100E),
				.b1(W2101E),
				.b2(W2102E),
				.b3(W2110E),
				.b4(W2111E),
				.b5(W2112E),
				.b6(W2120E),
				.b7(W2121E),
				.b8(W2122E),
				.c(c2E201)
);

ninexnine_unit ninexnine_unit_3219(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2100F),
				.b1(W2101F),
				.b2(W2102F),
				.b3(W2110F),
				.b4(W2111F),
				.b5(W2112F),
				.b6(W2120F),
				.b7(W2121F),
				.b8(W2122F),
				.c(c2F201)
);

assign C2201=c20201+c21201+c22201+c23201+c24201+c25201+c26201+c27201+c28201+c29201+c2A201+c2B201+c2C201+c2D201+c2E201+c2F201;
assign A2201=(C2201>=0)?1:0;

assign P3201=A2201;

ninexnine_unit ninexnine_unit_3220(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20211)
);

ninexnine_unit ninexnine_unit_3221(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21211)
);

ninexnine_unit ninexnine_unit_3222(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22211)
);

ninexnine_unit ninexnine_unit_3223(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23211)
);

ninexnine_unit ninexnine_unit_3224(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24211)
);

ninexnine_unit ninexnine_unit_3225(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25211)
);

ninexnine_unit ninexnine_unit_3226(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26211)
);

ninexnine_unit ninexnine_unit_3227(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27211)
);

ninexnine_unit ninexnine_unit_3228(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W21008),
				.b1(W21018),
				.b2(W21028),
				.b3(W21108),
				.b4(W21118),
				.b5(W21128),
				.b6(W21208),
				.b7(W21218),
				.b8(W21228),
				.c(c28211)
);

ninexnine_unit ninexnine_unit_3229(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W21009),
				.b1(W21019),
				.b2(W21029),
				.b3(W21109),
				.b4(W21119),
				.b5(W21129),
				.b6(W21209),
				.b7(W21219),
				.b8(W21229),
				.c(c29211)
);

ninexnine_unit ninexnine_unit_3230(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2100A),
				.b1(W2101A),
				.b2(W2102A),
				.b3(W2110A),
				.b4(W2111A),
				.b5(W2112A),
				.b6(W2120A),
				.b7(W2121A),
				.b8(W2122A),
				.c(c2A211)
);

ninexnine_unit ninexnine_unit_3231(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2100B),
				.b1(W2101B),
				.b2(W2102B),
				.b3(W2110B),
				.b4(W2111B),
				.b5(W2112B),
				.b6(W2120B),
				.b7(W2121B),
				.b8(W2122B),
				.c(c2B211)
);

ninexnine_unit ninexnine_unit_3232(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2100C),
				.b1(W2101C),
				.b2(W2102C),
				.b3(W2110C),
				.b4(W2111C),
				.b5(W2112C),
				.b6(W2120C),
				.b7(W2121C),
				.b8(W2122C),
				.c(c2C211)
);

ninexnine_unit ninexnine_unit_3233(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2100D),
				.b1(W2101D),
				.b2(W2102D),
				.b3(W2110D),
				.b4(W2111D),
				.b5(W2112D),
				.b6(W2120D),
				.b7(W2121D),
				.b8(W2122D),
				.c(c2D211)
);

ninexnine_unit ninexnine_unit_3234(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2100E),
				.b1(W2101E),
				.b2(W2102E),
				.b3(W2110E),
				.b4(W2111E),
				.b5(W2112E),
				.b6(W2120E),
				.b7(W2121E),
				.b8(W2122E),
				.c(c2E211)
);

ninexnine_unit ninexnine_unit_3235(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2100F),
				.b1(W2101F),
				.b2(W2102F),
				.b3(W2110F),
				.b4(W2111F),
				.b5(W2112F),
				.b6(W2120F),
				.b7(W2121F),
				.b8(W2122F),
				.c(c2F211)
);

assign C2211=c20211+c21211+c22211+c23211+c24211+c25211+c26211+c27211+c28211+c29211+c2A211+c2B211+c2C211+c2D211+c2E211+c2F211;
assign A2211=(C2211>=0)?1:0;

assign P3211=A2211;

ninexnine_unit ninexnine_unit_3236(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W21000),
				.b1(W21010),
				.b2(W21020),
				.b3(W21100),
				.b4(W21110),
				.b5(W21120),
				.b6(W21200),
				.b7(W21210),
				.b8(W21220),
				.c(c20221)
);

ninexnine_unit ninexnine_unit_3237(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W21001),
				.b1(W21011),
				.b2(W21021),
				.b3(W21101),
				.b4(W21111),
				.b5(W21121),
				.b6(W21201),
				.b7(W21211),
				.b8(W21221),
				.c(c21221)
);

ninexnine_unit ninexnine_unit_3238(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W21002),
				.b1(W21012),
				.b2(W21022),
				.b3(W21102),
				.b4(W21112),
				.b5(W21122),
				.b6(W21202),
				.b7(W21212),
				.b8(W21222),
				.c(c22221)
);

ninexnine_unit ninexnine_unit_3239(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W21003),
				.b1(W21013),
				.b2(W21023),
				.b3(W21103),
				.b4(W21113),
				.b5(W21123),
				.b6(W21203),
				.b7(W21213),
				.b8(W21223),
				.c(c23221)
);

ninexnine_unit ninexnine_unit_3240(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W21004),
				.b1(W21014),
				.b2(W21024),
				.b3(W21104),
				.b4(W21114),
				.b5(W21124),
				.b6(W21204),
				.b7(W21214),
				.b8(W21224),
				.c(c24221)
);

ninexnine_unit ninexnine_unit_3241(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W21005),
				.b1(W21015),
				.b2(W21025),
				.b3(W21105),
				.b4(W21115),
				.b5(W21125),
				.b6(W21205),
				.b7(W21215),
				.b8(W21225),
				.c(c25221)
);

ninexnine_unit ninexnine_unit_3242(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W21006),
				.b1(W21016),
				.b2(W21026),
				.b3(W21106),
				.b4(W21116),
				.b5(W21126),
				.b6(W21206),
				.b7(W21216),
				.b8(W21226),
				.c(c26221)
);

ninexnine_unit ninexnine_unit_3243(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W21007),
				.b1(W21017),
				.b2(W21027),
				.b3(W21107),
				.b4(W21117),
				.b5(W21127),
				.b6(W21207),
				.b7(W21217),
				.b8(W21227),
				.c(c27221)
);

ninexnine_unit ninexnine_unit_3244(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W21008),
				.b1(W21018),
				.b2(W21028),
				.b3(W21108),
				.b4(W21118),
				.b5(W21128),
				.b6(W21208),
				.b7(W21218),
				.b8(W21228),
				.c(c28221)
);

ninexnine_unit ninexnine_unit_3245(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W21009),
				.b1(W21019),
				.b2(W21029),
				.b3(W21109),
				.b4(W21119),
				.b5(W21129),
				.b6(W21209),
				.b7(W21219),
				.b8(W21229),
				.c(c29221)
);

ninexnine_unit ninexnine_unit_3246(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2100A),
				.b1(W2101A),
				.b2(W2102A),
				.b3(W2110A),
				.b4(W2111A),
				.b5(W2112A),
				.b6(W2120A),
				.b7(W2121A),
				.b8(W2122A),
				.c(c2A221)
);

ninexnine_unit ninexnine_unit_3247(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2100B),
				.b1(W2101B),
				.b2(W2102B),
				.b3(W2110B),
				.b4(W2111B),
				.b5(W2112B),
				.b6(W2120B),
				.b7(W2121B),
				.b8(W2122B),
				.c(c2B221)
);

ninexnine_unit ninexnine_unit_3248(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2100C),
				.b1(W2101C),
				.b2(W2102C),
				.b3(W2110C),
				.b4(W2111C),
				.b5(W2112C),
				.b6(W2120C),
				.b7(W2121C),
				.b8(W2122C),
				.c(c2C221)
);

ninexnine_unit ninexnine_unit_3249(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2100D),
				.b1(W2101D),
				.b2(W2102D),
				.b3(W2110D),
				.b4(W2111D),
				.b5(W2112D),
				.b6(W2120D),
				.b7(W2121D),
				.b8(W2122D),
				.c(c2D221)
);

ninexnine_unit ninexnine_unit_3250(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2100E),
				.b1(W2101E),
				.b2(W2102E),
				.b3(W2110E),
				.b4(W2111E),
				.b5(W2112E),
				.b6(W2120E),
				.b7(W2121E),
				.b8(W2122E),
				.c(c2E221)
);

ninexnine_unit ninexnine_unit_3251(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2100F),
				.b1(W2101F),
				.b2(W2102F),
				.b3(W2110F),
				.b4(W2111F),
				.b5(W2112F),
				.b6(W2120F),
				.b7(W2121F),
				.b8(W2122F),
				.c(c2F221)
);

assign C2221=c20221+c21221+c22221+c23221+c24221+c25221+c26221+c27221+c28221+c29221+c2A221+c2B221+c2C221+c2D221+c2E221+c2F221;
assign A2221=(C2221>=0)?1:0;

assign P3221=A2221;

ninexnine_unit ninexnine_unit_3252(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20002)
);

ninexnine_unit ninexnine_unit_3253(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21002)
);

ninexnine_unit ninexnine_unit_3254(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22002)
);

ninexnine_unit ninexnine_unit_3255(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23002)
);

ninexnine_unit ninexnine_unit_3256(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24002)
);

ninexnine_unit ninexnine_unit_3257(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25002)
);

ninexnine_unit ninexnine_unit_3258(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26002)
);

ninexnine_unit ninexnine_unit_3259(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27002)
);

ninexnine_unit ninexnine_unit_3260(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W22008),
				.b1(W22018),
				.b2(W22028),
				.b3(W22108),
				.b4(W22118),
				.b5(W22128),
				.b6(W22208),
				.b7(W22218),
				.b8(W22228),
				.c(c28002)
);

ninexnine_unit ninexnine_unit_3261(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W22009),
				.b1(W22019),
				.b2(W22029),
				.b3(W22109),
				.b4(W22119),
				.b5(W22129),
				.b6(W22209),
				.b7(W22219),
				.b8(W22229),
				.c(c29002)
);

ninexnine_unit ninexnine_unit_3262(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2200A),
				.b1(W2201A),
				.b2(W2202A),
				.b3(W2210A),
				.b4(W2211A),
				.b5(W2212A),
				.b6(W2220A),
				.b7(W2221A),
				.b8(W2222A),
				.c(c2A002)
);

ninexnine_unit ninexnine_unit_3263(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2200B),
				.b1(W2201B),
				.b2(W2202B),
				.b3(W2210B),
				.b4(W2211B),
				.b5(W2212B),
				.b6(W2220B),
				.b7(W2221B),
				.b8(W2222B),
				.c(c2B002)
);

ninexnine_unit ninexnine_unit_3264(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2200C),
				.b1(W2201C),
				.b2(W2202C),
				.b3(W2210C),
				.b4(W2211C),
				.b5(W2212C),
				.b6(W2220C),
				.b7(W2221C),
				.b8(W2222C),
				.c(c2C002)
);

ninexnine_unit ninexnine_unit_3265(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2200D),
				.b1(W2201D),
				.b2(W2202D),
				.b3(W2210D),
				.b4(W2211D),
				.b5(W2212D),
				.b6(W2220D),
				.b7(W2221D),
				.b8(W2222D),
				.c(c2D002)
);

ninexnine_unit ninexnine_unit_3266(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2200E),
				.b1(W2201E),
				.b2(W2202E),
				.b3(W2210E),
				.b4(W2211E),
				.b5(W2212E),
				.b6(W2220E),
				.b7(W2221E),
				.b8(W2222E),
				.c(c2E002)
);

ninexnine_unit ninexnine_unit_3267(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2200F),
				.b1(W2201F),
				.b2(W2202F),
				.b3(W2210F),
				.b4(W2211F),
				.b5(W2212F),
				.b6(W2220F),
				.b7(W2221F),
				.b8(W2222F),
				.c(c2F002)
);

assign C2002=c20002+c21002+c22002+c23002+c24002+c25002+c26002+c27002+c28002+c29002+c2A002+c2B002+c2C002+c2D002+c2E002+c2F002;
assign A2002=(C2002>=0)?1:0;

assign P3002=A2002;

ninexnine_unit ninexnine_unit_3268(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20012)
);

ninexnine_unit ninexnine_unit_3269(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21012)
);

ninexnine_unit ninexnine_unit_3270(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22012)
);

ninexnine_unit ninexnine_unit_3271(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23012)
);

ninexnine_unit ninexnine_unit_3272(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24012)
);

ninexnine_unit ninexnine_unit_3273(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25012)
);

ninexnine_unit ninexnine_unit_3274(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26012)
);

ninexnine_unit ninexnine_unit_3275(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27012)
);

ninexnine_unit ninexnine_unit_3276(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W22008),
				.b1(W22018),
				.b2(W22028),
				.b3(W22108),
				.b4(W22118),
				.b5(W22128),
				.b6(W22208),
				.b7(W22218),
				.b8(W22228),
				.c(c28012)
);

ninexnine_unit ninexnine_unit_3277(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W22009),
				.b1(W22019),
				.b2(W22029),
				.b3(W22109),
				.b4(W22119),
				.b5(W22129),
				.b6(W22209),
				.b7(W22219),
				.b8(W22229),
				.c(c29012)
);

ninexnine_unit ninexnine_unit_3278(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2200A),
				.b1(W2201A),
				.b2(W2202A),
				.b3(W2210A),
				.b4(W2211A),
				.b5(W2212A),
				.b6(W2220A),
				.b7(W2221A),
				.b8(W2222A),
				.c(c2A012)
);

ninexnine_unit ninexnine_unit_3279(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2200B),
				.b1(W2201B),
				.b2(W2202B),
				.b3(W2210B),
				.b4(W2211B),
				.b5(W2212B),
				.b6(W2220B),
				.b7(W2221B),
				.b8(W2222B),
				.c(c2B012)
);

ninexnine_unit ninexnine_unit_3280(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2200C),
				.b1(W2201C),
				.b2(W2202C),
				.b3(W2210C),
				.b4(W2211C),
				.b5(W2212C),
				.b6(W2220C),
				.b7(W2221C),
				.b8(W2222C),
				.c(c2C012)
);

ninexnine_unit ninexnine_unit_3281(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2200D),
				.b1(W2201D),
				.b2(W2202D),
				.b3(W2210D),
				.b4(W2211D),
				.b5(W2212D),
				.b6(W2220D),
				.b7(W2221D),
				.b8(W2222D),
				.c(c2D012)
);

ninexnine_unit ninexnine_unit_3282(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2200E),
				.b1(W2201E),
				.b2(W2202E),
				.b3(W2210E),
				.b4(W2211E),
				.b5(W2212E),
				.b6(W2220E),
				.b7(W2221E),
				.b8(W2222E),
				.c(c2E012)
);

ninexnine_unit ninexnine_unit_3283(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2200F),
				.b1(W2201F),
				.b2(W2202F),
				.b3(W2210F),
				.b4(W2211F),
				.b5(W2212F),
				.b6(W2220F),
				.b7(W2221F),
				.b8(W2222F),
				.c(c2F012)
);

assign C2012=c20012+c21012+c22012+c23012+c24012+c25012+c26012+c27012+c28012+c29012+c2A012+c2B012+c2C012+c2D012+c2E012+c2F012;
assign A2012=(C2012>=0)?1:0;

assign P3012=A2012;

ninexnine_unit ninexnine_unit_3284(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20022)
);

ninexnine_unit ninexnine_unit_3285(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21022)
);

ninexnine_unit ninexnine_unit_3286(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22022)
);

ninexnine_unit ninexnine_unit_3287(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23022)
);

ninexnine_unit ninexnine_unit_3288(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24022)
);

ninexnine_unit ninexnine_unit_3289(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25022)
);

ninexnine_unit ninexnine_unit_3290(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26022)
);

ninexnine_unit ninexnine_unit_3291(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27022)
);

ninexnine_unit ninexnine_unit_3292(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W22008),
				.b1(W22018),
				.b2(W22028),
				.b3(W22108),
				.b4(W22118),
				.b5(W22128),
				.b6(W22208),
				.b7(W22218),
				.b8(W22228),
				.c(c28022)
);

ninexnine_unit ninexnine_unit_3293(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W22009),
				.b1(W22019),
				.b2(W22029),
				.b3(W22109),
				.b4(W22119),
				.b5(W22129),
				.b6(W22209),
				.b7(W22219),
				.b8(W22229),
				.c(c29022)
);

ninexnine_unit ninexnine_unit_3294(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2200A),
				.b1(W2201A),
				.b2(W2202A),
				.b3(W2210A),
				.b4(W2211A),
				.b5(W2212A),
				.b6(W2220A),
				.b7(W2221A),
				.b8(W2222A),
				.c(c2A022)
);

ninexnine_unit ninexnine_unit_3295(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2200B),
				.b1(W2201B),
				.b2(W2202B),
				.b3(W2210B),
				.b4(W2211B),
				.b5(W2212B),
				.b6(W2220B),
				.b7(W2221B),
				.b8(W2222B),
				.c(c2B022)
);

ninexnine_unit ninexnine_unit_3296(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2200C),
				.b1(W2201C),
				.b2(W2202C),
				.b3(W2210C),
				.b4(W2211C),
				.b5(W2212C),
				.b6(W2220C),
				.b7(W2221C),
				.b8(W2222C),
				.c(c2C022)
);

ninexnine_unit ninexnine_unit_3297(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2200D),
				.b1(W2201D),
				.b2(W2202D),
				.b3(W2210D),
				.b4(W2211D),
				.b5(W2212D),
				.b6(W2220D),
				.b7(W2221D),
				.b8(W2222D),
				.c(c2D022)
);

ninexnine_unit ninexnine_unit_3298(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2200E),
				.b1(W2201E),
				.b2(W2202E),
				.b3(W2210E),
				.b4(W2211E),
				.b5(W2212E),
				.b6(W2220E),
				.b7(W2221E),
				.b8(W2222E),
				.c(c2E022)
);

ninexnine_unit ninexnine_unit_3299(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2200F),
				.b1(W2201F),
				.b2(W2202F),
				.b3(W2210F),
				.b4(W2211F),
				.b5(W2212F),
				.b6(W2220F),
				.b7(W2221F),
				.b8(W2222F),
				.c(c2F022)
);

assign C2022=c20022+c21022+c22022+c23022+c24022+c25022+c26022+c27022+c28022+c29022+c2A022+c2B022+c2C022+c2D022+c2E022+c2F022;
assign A2022=(C2022>=0)?1:0;

assign P3022=A2022;

ninexnine_unit ninexnine_unit_3300(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20102)
);

ninexnine_unit ninexnine_unit_3301(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21102)
);

ninexnine_unit ninexnine_unit_3302(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22102)
);

ninexnine_unit ninexnine_unit_3303(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23102)
);

ninexnine_unit ninexnine_unit_3304(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24102)
);

ninexnine_unit ninexnine_unit_3305(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25102)
);

ninexnine_unit ninexnine_unit_3306(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26102)
);

ninexnine_unit ninexnine_unit_3307(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27102)
);

ninexnine_unit ninexnine_unit_3308(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W22008),
				.b1(W22018),
				.b2(W22028),
				.b3(W22108),
				.b4(W22118),
				.b5(W22128),
				.b6(W22208),
				.b7(W22218),
				.b8(W22228),
				.c(c28102)
);

ninexnine_unit ninexnine_unit_3309(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W22009),
				.b1(W22019),
				.b2(W22029),
				.b3(W22109),
				.b4(W22119),
				.b5(W22129),
				.b6(W22209),
				.b7(W22219),
				.b8(W22229),
				.c(c29102)
);

ninexnine_unit ninexnine_unit_3310(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2200A),
				.b1(W2201A),
				.b2(W2202A),
				.b3(W2210A),
				.b4(W2211A),
				.b5(W2212A),
				.b6(W2220A),
				.b7(W2221A),
				.b8(W2222A),
				.c(c2A102)
);

ninexnine_unit ninexnine_unit_3311(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2200B),
				.b1(W2201B),
				.b2(W2202B),
				.b3(W2210B),
				.b4(W2211B),
				.b5(W2212B),
				.b6(W2220B),
				.b7(W2221B),
				.b8(W2222B),
				.c(c2B102)
);

ninexnine_unit ninexnine_unit_3312(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2200C),
				.b1(W2201C),
				.b2(W2202C),
				.b3(W2210C),
				.b4(W2211C),
				.b5(W2212C),
				.b6(W2220C),
				.b7(W2221C),
				.b8(W2222C),
				.c(c2C102)
);

ninexnine_unit ninexnine_unit_3313(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2200D),
				.b1(W2201D),
				.b2(W2202D),
				.b3(W2210D),
				.b4(W2211D),
				.b5(W2212D),
				.b6(W2220D),
				.b7(W2221D),
				.b8(W2222D),
				.c(c2D102)
);

ninexnine_unit ninexnine_unit_3314(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2200E),
				.b1(W2201E),
				.b2(W2202E),
				.b3(W2210E),
				.b4(W2211E),
				.b5(W2212E),
				.b6(W2220E),
				.b7(W2221E),
				.b8(W2222E),
				.c(c2E102)
);

ninexnine_unit ninexnine_unit_3315(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2200F),
				.b1(W2201F),
				.b2(W2202F),
				.b3(W2210F),
				.b4(W2211F),
				.b5(W2212F),
				.b6(W2220F),
				.b7(W2221F),
				.b8(W2222F),
				.c(c2F102)
);

assign C2102=c20102+c21102+c22102+c23102+c24102+c25102+c26102+c27102+c28102+c29102+c2A102+c2B102+c2C102+c2D102+c2E102+c2F102;
assign A2102=(C2102>=0)?1:0;

assign P3102=A2102;

ninexnine_unit ninexnine_unit_3316(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20112)
);

ninexnine_unit ninexnine_unit_3317(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21112)
);

ninexnine_unit ninexnine_unit_3318(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22112)
);

ninexnine_unit ninexnine_unit_3319(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23112)
);

ninexnine_unit ninexnine_unit_3320(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24112)
);

ninexnine_unit ninexnine_unit_3321(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25112)
);

ninexnine_unit ninexnine_unit_3322(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26112)
);

ninexnine_unit ninexnine_unit_3323(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27112)
);

ninexnine_unit ninexnine_unit_3324(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W22008),
				.b1(W22018),
				.b2(W22028),
				.b3(W22108),
				.b4(W22118),
				.b5(W22128),
				.b6(W22208),
				.b7(W22218),
				.b8(W22228),
				.c(c28112)
);

ninexnine_unit ninexnine_unit_3325(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W22009),
				.b1(W22019),
				.b2(W22029),
				.b3(W22109),
				.b4(W22119),
				.b5(W22129),
				.b6(W22209),
				.b7(W22219),
				.b8(W22229),
				.c(c29112)
);

ninexnine_unit ninexnine_unit_3326(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2200A),
				.b1(W2201A),
				.b2(W2202A),
				.b3(W2210A),
				.b4(W2211A),
				.b5(W2212A),
				.b6(W2220A),
				.b7(W2221A),
				.b8(W2222A),
				.c(c2A112)
);

ninexnine_unit ninexnine_unit_3327(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2200B),
				.b1(W2201B),
				.b2(W2202B),
				.b3(W2210B),
				.b4(W2211B),
				.b5(W2212B),
				.b6(W2220B),
				.b7(W2221B),
				.b8(W2222B),
				.c(c2B112)
);

ninexnine_unit ninexnine_unit_3328(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2200C),
				.b1(W2201C),
				.b2(W2202C),
				.b3(W2210C),
				.b4(W2211C),
				.b5(W2212C),
				.b6(W2220C),
				.b7(W2221C),
				.b8(W2222C),
				.c(c2C112)
);

ninexnine_unit ninexnine_unit_3329(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2200D),
				.b1(W2201D),
				.b2(W2202D),
				.b3(W2210D),
				.b4(W2211D),
				.b5(W2212D),
				.b6(W2220D),
				.b7(W2221D),
				.b8(W2222D),
				.c(c2D112)
);

ninexnine_unit ninexnine_unit_3330(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2200E),
				.b1(W2201E),
				.b2(W2202E),
				.b3(W2210E),
				.b4(W2211E),
				.b5(W2212E),
				.b6(W2220E),
				.b7(W2221E),
				.b8(W2222E),
				.c(c2E112)
);

ninexnine_unit ninexnine_unit_3331(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2200F),
				.b1(W2201F),
				.b2(W2202F),
				.b3(W2210F),
				.b4(W2211F),
				.b5(W2212F),
				.b6(W2220F),
				.b7(W2221F),
				.b8(W2222F),
				.c(c2F112)
);

assign C2112=c20112+c21112+c22112+c23112+c24112+c25112+c26112+c27112+c28112+c29112+c2A112+c2B112+c2C112+c2D112+c2E112+c2F112;
assign A2112=(C2112>=0)?1:0;

assign P3112=A2112;

ninexnine_unit ninexnine_unit_3332(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20122)
);

ninexnine_unit ninexnine_unit_3333(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21122)
);

ninexnine_unit ninexnine_unit_3334(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22122)
);

ninexnine_unit ninexnine_unit_3335(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23122)
);

ninexnine_unit ninexnine_unit_3336(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24122)
);

ninexnine_unit ninexnine_unit_3337(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25122)
);

ninexnine_unit ninexnine_unit_3338(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26122)
);

ninexnine_unit ninexnine_unit_3339(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27122)
);

ninexnine_unit ninexnine_unit_3340(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W22008),
				.b1(W22018),
				.b2(W22028),
				.b3(W22108),
				.b4(W22118),
				.b5(W22128),
				.b6(W22208),
				.b7(W22218),
				.b8(W22228),
				.c(c28122)
);

ninexnine_unit ninexnine_unit_3341(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W22009),
				.b1(W22019),
				.b2(W22029),
				.b3(W22109),
				.b4(W22119),
				.b5(W22129),
				.b6(W22209),
				.b7(W22219),
				.b8(W22229),
				.c(c29122)
);

ninexnine_unit ninexnine_unit_3342(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2200A),
				.b1(W2201A),
				.b2(W2202A),
				.b3(W2210A),
				.b4(W2211A),
				.b5(W2212A),
				.b6(W2220A),
				.b7(W2221A),
				.b8(W2222A),
				.c(c2A122)
);

ninexnine_unit ninexnine_unit_3343(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2200B),
				.b1(W2201B),
				.b2(W2202B),
				.b3(W2210B),
				.b4(W2211B),
				.b5(W2212B),
				.b6(W2220B),
				.b7(W2221B),
				.b8(W2222B),
				.c(c2B122)
);

ninexnine_unit ninexnine_unit_3344(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2200C),
				.b1(W2201C),
				.b2(W2202C),
				.b3(W2210C),
				.b4(W2211C),
				.b5(W2212C),
				.b6(W2220C),
				.b7(W2221C),
				.b8(W2222C),
				.c(c2C122)
);

ninexnine_unit ninexnine_unit_3345(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2200D),
				.b1(W2201D),
				.b2(W2202D),
				.b3(W2210D),
				.b4(W2211D),
				.b5(W2212D),
				.b6(W2220D),
				.b7(W2221D),
				.b8(W2222D),
				.c(c2D122)
);

ninexnine_unit ninexnine_unit_3346(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2200E),
				.b1(W2201E),
				.b2(W2202E),
				.b3(W2210E),
				.b4(W2211E),
				.b5(W2212E),
				.b6(W2220E),
				.b7(W2221E),
				.b8(W2222E),
				.c(c2E122)
);

ninexnine_unit ninexnine_unit_3347(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2200F),
				.b1(W2201F),
				.b2(W2202F),
				.b3(W2210F),
				.b4(W2211F),
				.b5(W2212F),
				.b6(W2220F),
				.b7(W2221F),
				.b8(W2222F),
				.c(c2F122)
);

assign C2122=c20122+c21122+c22122+c23122+c24122+c25122+c26122+c27122+c28122+c29122+c2A122+c2B122+c2C122+c2D122+c2E122+c2F122;
assign A2122=(C2122>=0)?1:0;

assign P3122=A2122;

ninexnine_unit ninexnine_unit_3348(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20202)
);

ninexnine_unit ninexnine_unit_3349(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21202)
);

ninexnine_unit ninexnine_unit_3350(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22202)
);

ninexnine_unit ninexnine_unit_3351(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23202)
);

ninexnine_unit ninexnine_unit_3352(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24202)
);

ninexnine_unit ninexnine_unit_3353(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25202)
);

ninexnine_unit ninexnine_unit_3354(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26202)
);

ninexnine_unit ninexnine_unit_3355(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27202)
);

ninexnine_unit ninexnine_unit_3356(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W22008),
				.b1(W22018),
				.b2(W22028),
				.b3(W22108),
				.b4(W22118),
				.b5(W22128),
				.b6(W22208),
				.b7(W22218),
				.b8(W22228),
				.c(c28202)
);

ninexnine_unit ninexnine_unit_3357(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W22009),
				.b1(W22019),
				.b2(W22029),
				.b3(W22109),
				.b4(W22119),
				.b5(W22129),
				.b6(W22209),
				.b7(W22219),
				.b8(W22229),
				.c(c29202)
);

ninexnine_unit ninexnine_unit_3358(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2200A),
				.b1(W2201A),
				.b2(W2202A),
				.b3(W2210A),
				.b4(W2211A),
				.b5(W2212A),
				.b6(W2220A),
				.b7(W2221A),
				.b8(W2222A),
				.c(c2A202)
);

ninexnine_unit ninexnine_unit_3359(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2200B),
				.b1(W2201B),
				.b2(W2202B),
				.b3(W2210B),
				.b4(W2211B),
				.b5(W2212B),
				.b6(W2220B),
				.b7(W2221B),
				.b8(W2222B),
				.c(c2B202)
);

ninexnine_unit ninexnine_unit_3360(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2200C),
				.b1(W2201C),
				.b2(W2202C),
				.b3(W2210C),
				.b4(W2211C),
				.b5(W2212C),
				.b6(W2220C),
				.b7(W2221C),
				.b8(W2222C),
				.c(c2C202)
);

ninexnine_unit ninexnine_unit_3361(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2200D),
				.b1(W2201D),
				.b2(W2202D),
				.b3(W2210D),
				.b4(W2211D),
				.b5(W2212D),
				.b6(W2220D),
				.b7(W2221D),
				.b8(W2222D),
				.c(c2D202)
);

ninexnine_unit ninexnine_unit_3362(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2200E),
				.b1(W2201E),
				.b2(W2202E),
				.b3(W2210E),
				.b4(W2211E),
				.b5(W2212E),
				.b6(W2220E),
				.b7(W2221E),
				.b8(W2222E),
				.c(c2E202)
);

ninexnine_unit ninexnine_unit_3363(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2200F),
				.b1(W2201F),
				.b2(W2202F),
				.b3(W2210F),
				.b4(W2211F),
				.b5(W2212F),
				.b6(W2220F),
				.b7(W2221F),
				.b8(W2222F),
				.c(c2F202)
);

assign C2202=c20202+c21202+c22202+c23202+c24202+c25202+c26202+c27202+c28202+c29202+c2A202+c2B202+c2C202+c2D202+c2E202+c2F202;
assign A2202=(C2202>=0)?1:0;

assign P3202=A2202;

ninexnine_unit ninexnine_unit_3364(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20212)
);

ninexnine_unit ninexnine_unit_3365(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21212)
);

ninexnine_unit ninexnine_unit_3366(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22212)
);

ninexnine_unit ninexnine_unit_3367(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23212)
);

ninexnine_unit ninexnine_unit_3368(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24212)
);

ninexnine_unit ninexnine_unit_3369(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25212)
);

ninexnine_unit ninexnine_unit_3370(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26212)
);

ninexnine_unit ninexnine_unit_3371(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27212)
);

ninexnine_unit ninexnine_unit_3372(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W22008),
				.b1(W22018),
				.b2(W22028),
				.b3(W22108),
				.b4(W22118),
				.b5(W22128),
				.b6(W22208),
				.b7(W22218),
				.b8(W22228),
				.c(c28212)
);

ninexnine_unit ninexnine_unit_3373(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W22009),
				.b1(W22019),
				.b2(W22029),
				.b3(W22109),
				.b4(W22119),
				.b5(W22129),
				.b6(W22209),
				.b7(W22219),
				.b8(W22229),
				.c(c29212)
);

ninexnine_unit ninexnine_unit_3374(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2200A),
				.b1(W2201A),
				.b2(W2202A),
				.b3(W2210A),
				.b4(W2211A),
				.b5(W2212A),
				.b6(W2220A),
				.b7(W2221A),
				.b8(W2222A),
				.c(c2A212)
);

ninexnine_unit ninexnine_unit_3375(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2200B),
				.b1(W2201B),
				.b2(W2202B),
				.b3(W2210B),
				.b4(W2211B),
				.b5(W2212B),
				.b6(W2220B),
				.b7(W2221B),
				.b8(W2222B),
				.c(c2B212)
);

ninexnine_unit ninexnine_unit_3376(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2200C),
				.b1(W2201C),
				.b2(W2202C),
				.b3(W2210C),
				.b4(W2211C),
				.b5(W2212C),
				.b6(W2220C),
				.b7(W2221C),
				.b8(W2222C),
				.c(c2C212)
);

ninexnine_unit ninexnine_unit_3377(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2200D),
				.b1(W2201D),
				.b2(W2202D),
				.b3(W2210D),
				.b4(W2211D),
				.b5(W2212D),
				.b6(W2220D),
				.b7(W2221D),
				.b8(W2222D),
				.c(c2D212)
);

ninexnine_unit ninexnine_unit_3378(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2200E),
				.b1(W2201E),
				.b2(W2202E),
				.b3(W2210E),
				.b4(W2211E),
				.b5(W2212E),
				.b6(W2220E),
				.b7(W2221E),
				.b8(W2222E),
				.c(c2E212)
);

ninexnine_unit ninexnine_unit_3379(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2200F),
				.b1(W2201F),
				.b2(W2202F),
				.b3(W2210F),
				.b4(W2211F),
				.b5(W2212F),
				.b6(W2220F),
				.b7(W2221F),
				.b8(W2222F),
				.c(c2F212)
);

assign C2212=c20212+c21212+c22212+c23212+c24212+c25212+c26212+c27212+c28212+c29212+c2A212+c2B212+c2C212+c2D212+c2E212+c2F212;
assign A2212=(C2212>=0)?1:0;

assign P3212=A2212;

ninexnine_unit ninexnine_unit_3380(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W22000),
				.b1(W22010),
				.b2(W22020),
				.b3(W22100),
				.b4(W22110),
				.b5(W22120),
				.b6(W22200),
				.b7(W22210),
				.b8(W22220),
				.c(c20222)
);

ninexnine_unit ninexnine_unit_3381(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W22001),
				.b1(W22011),
				.b2(W22021),
				.b3(W22101),
				.b4(W22111),
				.b5(W22121),
				.b6(W22201),
				.b7(W22211),
				.b8(W22221),
				.c(c21222)
);

ninexnine_unit ninexnine_unit_3382(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W22002),
				.b1(W22012),
				.b2(W22022),
				.b3(W22102),
				.b4(W22112),
				.b5(W22122),
				.b6(W22202),
				.b7(W22212),
				.b8(W22222),
				.c(c22222)
);

ninexnine_unit ninexnine_unit_3383(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W22003),
				.b1(W22013),
				.b2(W22023),
				.b3(W22103),
				.b4(W22113),
				.b5(W22123),
				.b6(W22203),
				.b7(W22213),
				.b8(W22223),
				.c(c23222)
);

ninexnine_unit ninexnine_unit_3384(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W22004),
				.b1(W22014),
				.b2(W22024),
				.b3(W22104),
				.b4(W22114),
				.b5(W22124),
				.b6(W22204),
				.b7(W22214),
				.b8(W22224),
				.c(c24222)
);

ninexnine_unit ninexnine_unit_3385(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W22005),
				.b1(W22015),
				.b2(W22025),
				.b3(W22105),
				.b4(W22115),
				.b5(W22125),
				.b6(W22205),
				.b7(W22215),
				.b8(W22225),
				.c(c25222)
);

ninexnine_unit ninexnine_unit_3386(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W22006),
				.b1(W22016),
				.b2(W22026),
				.b3(W22106),
				.b4(W22116),
				.b5(W22126),
				.b6(W22206),
				.b7(W22216),
				.b8(W22226),
				.c(c26222)
);

ninexnine_unit ninexnine_unit_3387(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W22007),
				.b1(W22017),
				.b2(W22027),
				.b3(W22107),
				.b4(W22117),
				.b5(W22127),
				.b6(W22207),
				.b7(W22217),
				.b8(W22227),
				.c(c27222)
);

ninexnine_unit ninexnine_unit_3388(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W22008),
				.b1(W22018),
				.b2(W22028),
				.b3(W22108),
				.b4(W22118),
				.b5(W22128),
				.b6(W22208),
				.b7(W22218),
				.b8(W22228),
				.c(c28222)
);

ninexnine_unit ninexnine_unit_3389(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W22009),
				.b1(W22019),
				.b2(W22029),
				.b3(W22109),
				.b4(W22119),
				.b5(W22129),
				.b6(W22209),
				.b7(W22219),
				.b8(W22229),
				.c(c29222)
);

ninexnine_unit ninexnine_unit_3390(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2200A),
				.b1(W2201A),
				.b2(W2202A),
				.b3(W2210A),
				.b4(W2211A),
				.b5(W2212A),
				.b6(W2220A),
				.b7(W2221A),
				.b8(W2222A),
				.c(c2A222)
);

ninexnine_unit ninexnine_unit_3391(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2200B),
				.b1(W2201B),
				.b2(W2202B),
				.b3(W2210B),
				.b4(W2211B),
				.b5(W2212B),
				.b6(W2220B),
				.b7(W2221B),
				.b8(W2222B),
				.c(c2B222)
);

ninexnine_unit ninexnine_unit_3392(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2200C),
				.b1(W2201C),
				.b2(W2202C),
				.b3(W2210C),
				.b4(W2211C),
				.b5(W2212C),
				.b6(W2220C),
				.b7(W2221C),
				.b8(W2222C),
				.c(c2C222)
);

ninexnine_unit ninexnine_unit_3393(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2200D),
				.b1(W2201D),
				.b2(W2202D),
				.b3(W2210D),
				.b4(W2211D),
				.b5(W2212D),
				.b6(W2220D),
				.b7(W2221D),
				.b8(W2222D),
				.c(c2D222)
);

ninexnine_unit ninexnine_unit_3394(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2200E),
				.b1(W2201E),
				.b2(W2202E),
				.b3(W2210E),
				.b4(W2211E),
				.b5(W2212E),
				.b6(W2220E),
				.b7(W2221E),
				.b8(W2222E),
				.c(c2E222)
);

ninexnine_unit ninexnine_unit_3395(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2200F),
				.b1(W2201F),
				.b2(W2202F),
				.b3(W2210F),
				.b4(W2211F),
				.b5(W2212F),
				.b6(W2220F),
				.b7(W2221F),
				.b8(W2222F),
				.c(c2F222)
);

assign C2222=c20222+c21222+c22222+c23222+c24222+c25222+c26222+c27222+c28222+c29222+c2A222+c2B222+c2C222+c2D222+c2E222+c2F222;
assign A2222=(C2222>=0)?1:0;

assign P3222=A2222;

ninexnine_unit ninexnine_unit_3396(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20003)
);

ninexnine_unit ninexnine_unit_3397(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21003)
);

ninexnine_unit ninexnine_unit_3398(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22003)
);

ninexnine_unit ninexnine_unit_3399(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23003)
);

ninexnine_unit ninexnine_unit_3400(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24003)
);

ninexnine_unit ninexnine_unit_3401(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25003)
);

ninexnine_unit ninexnine_unit_3402(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26003)
);

ninexnine_unit ninexnine_unit_3403(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27003)
);

ninexnine_unit ninexnine_unit_3404(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W23008),
				.b1(W23018),
				.b2(W23028),
				.b3(W23108),
				.b4(W23118),
				.b5(W23128),
				.b6(W23208),
				.b7(W23218),
				.b8(W23228),
				.c(c28003)
);

ninexnine_unit ninexnine_unit_3405(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W23009),
				.b1(W23019),
				.b2(W23029),
				.b3(W23109),
				.b4(W23119),
				.b5(W23129),
				.b6(W23209),
				.b7(W23219),
				.b8(W23229),
				.c(c29003)
);

ninexnine_unit ninexnine_unit_3406(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2300A),
				.b1(W2301A),
				.b2(W2302A),
				.b3(W2310A),
				.b4(W2311A),
				.b5(W2312A),
				.b6(W2320A),
				.b7(W2321A),
				.b8(W2322A),
				.c(c2A003)
);

ninexnine_unit ninexnine_unit_3407(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2300B),
				.b1(W2301B),
				.b2(W2302B),
				.b3(W2310B),
				.b4(W2311B),
				.b5(W2312B),
				.b6(W2320B),
				.b7(W2321B),
				.b8(W2322B),
				.c(c2B003)
);

ninexnine_unit ninexnine_unit_3408(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2300C),
				.b1(W2301C),
				.b2(W2302C),
				.b3(W2310C),
				.b4(W2311C),
				.b5(W2312C),
				.b6(W2320C),
				.b7(W2321C),
				.b8(W2322C),
				.c(c2C003)
);

ninexnine_unit ninexnine_unit_3409(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2300D),
				.b1(W2301D),
				.b2(W2302D),
				.b3(W2310D),
				.b4(W2311D),
				.b5(W2312D),
				.b6(W2320D),
				.b7(W2321D),
				.b8(W2322D),
				.c(c2D003)
);

ninexnine_unit ninexnine_unit_3410(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2300E),
				.b1(W2301E),
				.b2(W2302E),
				.b3(W2310E),
				.b4(W2311E),
				.b5(W2312E),
				.b6(W2320E),
				.b7(W2321E),
				.b8(W2322E),
				.c(c2E003)
);

ninexnine_unit ninexnine_unit_3411(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2300F),
				.b1(W2301F),
				.b2(W2302F),
				.b3(W2310F),
				.b4(W2311F),
				.b5(W2312F),
				.b6(W2320F),
				.b7(W2321F),
				.b8(W2322F),
				.c(c2F003)
);

assign C2003=c20003+c21003+c22003+c23003+c24003+c25003+c26003+c27003+c28003+c29003+c2A003+c2B003+c2C003+c2D003+c2E003+c2F003;
assign A2003=(C2003>=0)?1:0;

assign P3003=A2003;

ninexnine_unit ninexnine_unit_3412(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20013)
);

ninexnine_unit ninexnine_unit_3413(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21013)
);

ninexnine_unit ninexnine_unit_3414(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22013)
);

ninexnine_unit ninexnine_unit_3415(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23013)
);

ninexnine_unit ninexnine_unit_3416(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24013)
);

ninexnine_unit ninexnine_unit_3417(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25013)
);

ninexnine_unit ninexnine_unit_3418(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26013)
);

ninexnine_unit ninexnine_unit_3419(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27013)
);

ninexnine_unit ninexnine_unit_3420(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W23008),
				.b1(W23018),
				.b2(W23028),
				.b3(W23108),
				.b4(W23118),
				.b5(W23128),
				.b6(W23208),
				.b7(W23218),
				.b8(W23228),
				.c(c28013)
);

ninexnine_unit ninexnine_unit_3421(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W23009),
				.b1(W23019),
				.b2(W23029),
				.b3(W23109),
				.b4(W23119),
				.b5(W23129),
				.b6(W23209),
				.b7(W23219),
				.b8(W23229),
				.c(c29013)
);

ninexnine_unit ninexnine_unit_3422(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2300A),
				.b1(W2301A),
				.b2(W2302A),
				.b3(W2310A),
				.b4(W2311A),
				.b5(W2312A),
				.b6(W2320A),
				.b7(W2321A),
				.b8(W2322A),
				.c(c2A013)
);

ninexnine_unit ninexnine_unit_3423(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2300B),
				.b1(W2301B),
				.b2(W2302B),
				.b3(W2310B),
				.b4(W2311B),
				.b5(W2312B),
				.b6(W2320B),
				.b7(W2321B),
				.b8(W2322B),
				.c(c2B013)
);

ninexnine_unit ninexnine_unit_3424(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2300C),
				.b1(W2301C),
				.b2(W2302C),
				.b3(W2310C),
				.b4(W2311C),
				.b5(W2312C),
				.b6(W2320C),
				.b7(W2321C),
				.b8(W2322C),
				.c(c2C013)
);

ninexnine_unit ninexnine_unit_3425(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2300D),
				.b1(W2301D),
				.b2(W2302D),
				.b3(W2310D),
				.b4(W2311D),
				.b5(W2312D),
				.b6(W2320D),
				.b7(W2321D),
				.b8(W2322D),
				.c(c2D013)
);

ninexnine_unit ninexnine_unit_3426(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2300E),
				.b1(W2301E),
				.b2(W2302E),
				.b3(W2310E),
				.b4(W2311E),
				.b5(W2312E),
				.b6(W2320E),
				.b7(W2321E),
				.b8(W2322E),
				.c(c2E013)
);

ninexnine_unit ninexnine_unit_3427(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2300F),
				.b1(W2301F),
				.b2(W2302F),
				.b3(W2310F),
				.b4(W2311F),
				.b5(W2312F),
				.b6(W2320F),
				.b7(W2321F),
				.b8(W2322F),
				.c(c2F013)
);

assign C2013=c20013+c21013+c22013+c23013+c24013+c25013+c26013+c27013+c28013+c29013+c2A013+c2B013+c2C013+c2D013+c2E013+c2F013;
assign A2013=(C2013>=0)?1:0;

assign P3013=A2013;

ninexnine_unit ninexnine_unit_3428(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20023)
);

ninexnine_unit ninexnine_unit_3429(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21023)
);

ninexnine_unit ninexnine_unit_3430(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22023)
);

ninexnine_unit ninexnine_unit_3431(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23023)
);

ninexnine_unit ninexnine_unit_3432(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24023)
);

ninexnine_unit ninexnine_unit_3433(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25023)
);

ninexnine_unit ninexnine_unit_3434(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26023)
);

ninexnine_unit ninexnine_unit_3435(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27023)
);

ninexnine_unit ninexnine_unit_3436(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W23008),
				.b1(W23018),
				.b2(W23028),
				.b3(W23108),
				.b4(W23118),
				.b5(W23128),
				.b6(W23208),
				.b7(W23218),
				.b8(W23228),
				.c(c28023)
);

ninexnine_unit ninexnine_unit_3437(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W23009),
				.b1(W23019),
				.b2(W23029),
				.b3(W23109),
				.b4(W23119),
				.b5(W23129),
				.b6(W23209),
				.b7(W23219),
				.b8(W23229),
				.c(c29023)
);

ninexnine_unit ninexnine_unit_3438(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2300A),
				.b1(W2301A),
				.b2(W2302A),
				.b3(W2310A),
				.b4(W2311A),
				.b5(W2312A),
				.b6(W2320A),
				.b7(W2321A),
				.b8(W2322A),
				.c(c2A023)
);

ninexnine_unit ninexnine_unit_3439(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2300B),
				.b1(W2301B),
				.b2(W2302B),
				.b3(W2310B),
				.b4(W2311B),
				.b5(W2312B),
				.b6(W2320B),
				.b7(W2321B),
				.b8(W2322B),
				.c(c2B023)
);

ninexnine_unit ninexnine_unit_3440(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2300C),
				.b1(W2301C),
				.b2(W2302C),
				.b3(W2310C),
				.b4(W2311C),
				.b5(W2312C),
				.b6(W2320C),
				.b7(W2321C),
				.b8(W2322C),
				.c(c2C023)
);

ninexnine_unit ninexnine_unit_3441(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2300D),
				.b1(W2301D),
				.b2(W2302D),
				.b3(W2310D),
				.b4(W2311D),
				.b5(W2312D),
				.b6(W2320D),
				.b7(W2321D),
				.b8(W2322D),
				.c(c2D023)
);

ninexnine_unit ninexnine_unit_3442(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2300E),
				.b1(W2301E),
				.b2(W2302E),
				.b3(W2310E),
				.b4(W2311E),
				.b5(W2312E),
				.b6(W2320E),
				.b7(W2321E),
				.b8(W2322E),
				.c(c2E023)
);

ninexnine_unit ninexnine_unit_3443(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2300F),
				.b1(W2301F),
				.b2(W2302F),
				.b3(W2310F),
				.b4(W2311F),
				.b5(W2312F),
				.b6(W2320F),
				.b7(W2321F),
				.b8(W2322F),
				.c(c2F023)
);

assign C2023=c20023+c21023+c22023+c23023+c24023+c25023+c26023+c27023+c28023+c29023+c2A023+c2B023+c2C023+c2D023+c2E023+c2F023;
assign A2023=(C2023>=0)?1:0;

assign P3023=A2023;

ninexnine_unit ninexnine_unit_3444(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20103)
);

ninexnine_unit ninexnine_unit_3445(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21103)
);

ninexnine_unit ninexnine_unit_3446(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22103)
);

ninexnine_unit ninexnine_unit_3447(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23103)
);

ninexnine_unit ninexnine_unit_3448(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24103)
);

ninexnine_unit ninexnine_unit_3449(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25103)
);

ninexnine_unit ninexnine_unit_3450(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26103)
);

ninexnine_unit ninexnine_unit_3451(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27103)
);

ninexnine_unit ninexnine_unit_3452(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W23008),
				.b1(W23018),
				.b2(W23028),
				.b3(W23108),
				.b4(W23118),
				.b5(W23128),
				.b6(W23208),
				.b7(W23218),
				.b8(W23228),
				.c(c28103)
);

ninexnine_unit ninexnine_unit_3453(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W23009),
				.b1(W23019),
				.b2(W23029),
				.b3(W23109),
				.b4(W23119),
				.b5(W23129),
				.b6(W23209),
				.b7(W23219),
				.b8(W23229),
				.c(c29103)
);

ninexnine_unit ninexnine_unit_3454(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2300A),
				.b1(W2301A),
				.b2(W2302A),
				.b3(W2310A),
				.b4(W2311A),
				.b5(W2312A),
				.b6(W2320A),
				.b7(W2321A),
				.b8(W2322A),
				.c(c2A103)
);

ninexnine_unit ninexnine_unit_3455(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2300B),
				.b1(W2301B),
				.b2(W2302B),
				.b3(W2310B),
				.b4(W2311B),
				.b5(W2312B),
				.b6(W2320B),
				.b7(W2321B),
				.b8(W2322B),
				.c(c2B103)
);

ninexnine_unit ninexnine_unit_3456(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2300C),
				.b1(W2301C),
				.b2(W2302C),
				.b3(W2310C),
				.b4(W2311C),
				.b5(W2312C),
				.b6(W2320C),
				.b7(W2321C),
				.b8(W2322C),
				.c(c2C103)
);

ninexnine_unit ninexnine_unit_3457(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2300D),
				.b1(W2301D),
				.b2(W2302D),
				.b3(W2310D),
				.b4(W2311D),
				.b5(W2312D),
				.b6(W2320D),
				.b7(W2321D),
				.b8(W2322D),
				.c(c2D103)
);

ninexnine_unit ninexnine_unit_3458(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2300E),
				.b1(W2301E),
				.b2(W2302E),
				.b3(W2310E),
				.b4(W2311E),
				.b5(W2312E),
				.b6(W2320E),
				.b7(W2321E),
				.b8(W2322E),
				.c(c2E103)
);

ninexnine_unit ninexnine_unit_3459(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2300F),
				.b1(W2301F),
				.b2(W2302F),
				.b3(W2310F),
				.b4(W2311F),
				.b5(W2312F),
				.b6(W2320F),
				.b7(W2321F),
				.b8(W2322F),
				.c(c2F103)
);

assign C2103=c20103+c21103+c22103+c23103+c24103+c25103+c26103+c27103+c28103+c29103+c2A103+c2B103+c2C103+c2D103+c2E103+c2F103;
assign A2103=(C2103>=0)?1:0;

assign P3103=A2103;

ninexnine_unit ninexnine_unit_3460(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20113)
);

ninexnine_unit ninexnine_unit_3461(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21113)
);

ninexnine_unit ninexnine_unit_3462(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22113)
);

ninexnine_unit ninexnine_unit_3463(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23113)
);

ninexnine_unit ninexnine_unit_3464(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24113)
);

ninexnine_unit ninexnine_unit_3465(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25113)
);

ninexnine_unit ninexnine_unit_3466(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26113)
);

ninexnine_unit ninexnine_unit_3467(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27113)
);

ninexnine_unit ninexnine_unit_3468(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W23008),
				.b1(W23018),
				.b2(W23028),
				.b3(W23108),
				.b4(W23118),
				.b5(W23128),
				.b6(W23208),
				.b7(W23218),
				.b8(W23228),
				.c(c28113)
);

ninexnine_unit ninexnine_unit_3469(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W23009),
				.b1(W23019),
				.b2(W23029),
				.b3(W23109),
				.b4(W23119),
				.b5(W23129),
				.b6(W23209),
				.b7(W23219),
				.b8(W23229),
				.c(c29113)
);

ninexnine_unit ninexnine_unit_3470(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2300A),
				.b1(W2301A),
				.b2(W2302A),
				.b3(W2310A),
				.b4(W2311A),
				.b5(W2312A),
				.b6(W2320A),
				.b7(W2321A),
				.b8(W2322A),
				.c(c2A113)
);

ninexnine_unit ninexnine_unit_3471(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2300B),
				.b1(W2301B),
				.b2(W2302B),
				.b3(W2310B),
				.b4(W2311B),
				.b5(W2312B),
				.b6(W2320B),
				.b7(W2321B),
				.b8(W2322B),
				.c(c2B113)
);

ninexnine_unit ninexnine_unit_3472(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2300C),
				.b1(W2301C),
				.b2(W2302C),
				.b3(W2310C),
				.b4(W2311C),
				.b5(W2312C),
				.b6(W2320C),
				.b7(W2321C),
				.b8(W2322C),
				.c(c2C113)
);

ninexnine_unit ninexnine_unit_3473(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2300D),
				.b1(W2301D),
				.b2(W2302D),
				.b3(W2310D),
				.b4(W2311D),
				.b5(W2312D),
				.b6(W2320D),
				.b7(W2321D),
				.b8(W2322D),
				.c(c2D113)
);

ninexnine_unit ninexnine_unit_3474(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2300E),
				.b1(W2301E),
				.b2(W2302E),
				.b3(W2310E),
				.b4(W2311E),
				.b5(W2312E),
				.b6(W2320E),
				.b7(W2321E),
				.b8(W2322E),
				.c(c2E113)
);

ninexnine_unit ninexnine_unit_3475(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2300F),
				.b1(W2301F),
				.b2(W2302F),
				.b3(W2310F),
				.b4(W2311F),
				.b5(W2312F),
				.b6(W2320F),
				.b7(W2321F),
				.b8(W2322F),
				.c(c2F113)
);

assign C2113=c20113+c21113+c22113+c23113+c24113+c25113+c26113+c27113+c28113+c29113+c2A113+c2B113+c2C113+c2D113+c2E113+c2F113;
assign A2113=(C2113>=0)?1:0;

assign P3113=A2113;

ninexnine_unit ninexnine_unit_3476(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20123)
);

ninexnine_unit ninexnine_unit_3477(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21123)
);

ninexnine_unit ninexnine_unit_3478(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22123)
);

ninexnine_unit ninexnine_unit_3479(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23123)
);

ninexnine_unit ninexnine_unit_3480(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24123)
);

ninexnine_unit ninexnine_unit_3481(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25123)
);

ninexnine_unit ninexnine_unit_3482(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26123)
);

ninexnine_unit ninexnine_unit_3483(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27123)
);

ninexnine_unit ninexnine_unit_3484(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W23008),
				.b1(W23018),
				.b2(W23028),
				.b3(W23108),
				.b4(W23118),
				.b5(W23128),
				.b6(W23208),
				.b7(W23218),
				.b8(W23228),
				.c(c28123)
);

ninexnine_unit ninexnine_unit_3485(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W23009),
				.b1(W23019),
				.b2(W23029),
				.b3(W23109),
				.b4(W23119),
				.b5(W23129),
				.b6(W23209),
				.b7(W23219),
				.b8(W23229),
				.c(c29123)
);

ninexnine_unit ninexnine_unit_3486(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2300A),
				.b1(W2301A),
				.b2(W2302A),
				.b3(W2310A),
				.b4(W2311A),
				.b5(W2312A),
				.b6(W2320A),
				.b7(W2321A),
				.b8(W2322A),
				.c(c2A123)
);

ninexnine_unit ninexnine_unit_3487(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2300B),
				.b1(W2301B),
				.b2(W2302B),
				.b3(W2310B),
				.b4(W2311B),
				.b5(W2312B),
				.b6(W2320B),
				.b7(W2321B),
				.b8(W2322B),
				.c(c2B123)
);

ninexnine_unit ninexnine_unit_3488(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2300C),
				.b1(W2301C),
				.b2(W2302C),
				.b3(W2310C),
				.b4(W2311C),
				.b5(W2312C),
				.b6(W2320C),
				.b7(W2321C),
				.b8(W2322C),
				.c(c2C123)
);

ninexnine_unit ninexnine_unit_3489(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2300D),
				.b1(W2301D),
				.b2(W2302D),
				.b3(W2310D),
				.b4(W2311D),
				.b5(W2312D),
				.b6(W2320D),
				.b7(W2321D),
				.b8(W2322D),
				.c(c2D123)
);

ninexnine_unit ninexnine_unit_3490(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2300E),
				.b1(W2301E),
				.b2(W2302E),
				.b3(W2310E),
				.b4(W2311E),
				.b5(W2312E),
				.b6(W2320E),
				.b7(W2321E),
				.b8(W2322E),
				.c(c2E123)
);

ninexnine_unit ninexnine_unit_3491(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2300F),
				.b1(W2301F),
				.b2(W2302F),
				.b3(W2310F),
				.b4(W2311F),
				.b5(W2312F),
				.b6(W2320F),
				.b7(W2321F),
				.b8(W2322F),
				.c(c2F123)
);

assign C2123=c20123+c21123+c22123+c23123+c24123+c25123+c26123+c27123+c28123+c29123+c2A123+c2B123+c2C123+c2D123+c2E123+c2F123;
assign A2123=(C2123>=0)?1:0;

assign P3123=A2123;

ninexnine_unit ninexnine_unit_3492(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20203)
);

ninexnine_unit ninexnine_unit_3493(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21203)
);

ninexnine_unit ninexnine_unit_3494(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22203)
);

ninexnine_unit ninexnine_unit_3495(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23203)
);

ninexnine_unit ninexnine_unit_3496(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24203)
);

ninexnine_unit ninexnine_unit_3497(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25203)
);

ninexnine_unit ninexnine_unit_3498(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26203)
);

ninexnine_unit ninexnine_unit_3499(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27203)
);

ninexnine_unit ninexnine_unit_3500(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W23008),
				.b1(W23018),
				.b2(W23028),
				.b3(W23108),
				.b4(W23118),
				.b5(W23128),
				.b6(W23208),
				.b7(W23218),
				.b8(W23228),
				.c(c28203)
);

ninexnine_unit ninexnine_unit_3501(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W23009),
				.b1(W23019),
				.b2(W23029),
				.b3(W23109),
				.b4(W23119),
				.b5(W23129),
				.b6(W23209),
				.b7(W23219),
				.b8(W23229),
				.c(c29203)
);

ninexnine_unit ninexnine_unit_3502(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2300A),
				.b1(W2301A),
				.b2(W2302A),
				.b3(W2310A),
				.b4(W2311A),
				.b5(W2312A),
				.b6(W2320A),
				.b7(W2321A),
				.b8(W2322A),
				.c(c2A203)
);

ninexnine_unit ninexnine_unit_3503(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2300B),
				.b1(W2301B),
				.b2(W2302B),
				.b3(W2310B),
				.b4(W2311B),
				.b5(W2312B),
				.b6(W2320B),
				.b7(W2321B),
				.b8(W2322B),
				.c(c2B203)
);

ninexnine_unit ninexnine_unit_3504(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2300C),
				.b1(W2301C),
				.b2(W2302C),
				.b3(W2310C),
				.b4(W2311C),
				.b5(W2312C),
				.b6(W2320C),
				.b7(W2321C),
				.b8(W2322C),
				.c(c2C203)
);

ninexnine_unit ninexnine_unit_3505(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2300D),
				.b1(W2301D),
				.b2(W2302D),
				.b3(W2310D),
				.b4(W2311D),
				.b5(W2312D),
				.b6(W2320D),
				.b7(W2321D),
				.b8(W2322D),
				.c(c2D203)
);

ninexnine_unit ninexnine_unit_3506(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2300E),
				.b1(W2301E),
				.b2(W2302E),
				.b3(W2310E),
				.b4(W2311E),
				.b5(W2312E),
				.b6(W2320E),
				.b7(W2321E),
				.b8(W2322E),
				.c(c2E203)
);

ninexnine_unit ninexnine_unit_3507(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2300F),
				.b1(W2301F),
				.b2(W2302F),
				.b3(W2310F),
				.b4(W2311F),
				.b5(W2312F),
				.b6(W2320F),
				.b7(W2321F),
				.b8(W2322F),
				.c(c2F203)
);

assign C2203=c20203+c21203+c22203+c23203+c24203+c25203+c26203+c27203+c28203+c29203+c2A203+c2B203+c2C203+c2D203+c2E203+c2F203;
assign A2203=(C2203>=0)?1:0;

assign P3203=A2203;

ninexnine_unit ninexnine_unit_3508(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20213)
);

ninexnine_unit ninexnine_unit_3509(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21213)
);

ninexnine_unit ninexnine_unit_3510(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22213)
);

ninexnine_unit ninexnine_unit_3511(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23213)
);

ninexnine_unit ninexnine_unit_3512(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24213)
);

ninexnine_unit ninexnine_unit_3513(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25213)
);

ninexnine_unit ninexnine_unit_3514(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26213)
);

ninexnine_unit ninexnine_unit_3515(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27213)
);

ninexnine_unit ninexnine_unit_3516(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W23008),
				.b1(W23018),
				.b2(W23028),
				.b3(W23108),
				.b4(W23118),
				.b5(W23128),
				.b6(W23208),
				.b7(W23218),
				.b8(W23228),
				.c(c28213)
);

ninexnine_unit ninexnine_unit_3517(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W23009),
				.b1(W23019),
				.b2(W23029),
				.b3(W23109),
				.b4(W23119),
				.b5(W23129),
				.b6(W23209),
				.b7(W23219),
				.b8(W23229),
				.c(c29213)
);

ninexnine_unit ninexnine_unit_3518(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2300A),
				.b1(W2301A),
				.b2(W2302A),
				.b3(W2310A),
				.b4(W2311A),
				.b5(W2312A),
				.b6(W2320A),
				.b7(W2321A),
				.b8(W2322A),
				.c(c2A213)
);

ninexnine_unit ninexnine_unit_3519(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2300B),
				.b1(W2301B),
				.b2(W2302B),
				.b3(W2310B),
				.b4(W2311B),
				.b5(W2312B),
				.b6(W2320B),
				.b7(W2321B),
				.b8(W2322B),
				.c(c2B213)
);

ninexnine_unit ninexnine_unit_3520(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2300C),
				.b1(W2301C),
				.b2(W2302C),
				.b3(W2310C),
				.b4(W2311C),
				.b5(W2312C),
				.b6(W2320C),
				.b7(W2321C),
				.b8(W2322C),
				.c(c2C213)
);

ninexnine_unit ninexnine_unit_3521(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2300D),
				.b1(W2301D),
				.b2(W2302D),
				.b3(W2310D),
				.b4(W2311D),
				.b5(W2312D),
				.b6(W2320D),
				.b7(W2321D),
				.b8(W2322D),
				.c(c2D213)
);

ninexnine_unit ninexnine_unit_3522(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2300E),
				.b1(W2301E),
				.b2(W2302E),
				.b3(W2310E),
				.b4(W2311E),
				.b5(W2312E),
				.b6(W2320E),
				.b7(W2321E),
				.b8(W2322E),
				.c(c2E213)
);

ninexnine_unit ninexnine_unit_3523(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2300F),
				.b1(W2301F),
				.b2(W2302F),
				.b3(W2310F),
				.b4(W2311F),
				.b5(W2312F),
				.b6(W2320F),
				.b7(W2321F),
				.b8(W2322F),
				.c(c2F213)
);

assign C2213=c20213+c21213+c22213+c23213+c24213+c25213+c26213+c27213+c28213+c29213+c2A213+c2B213+c2C213+c2D213+c2E213+c2F213;
assign A2213=(C2213>=0)?1:0;

assign P3213=A2213;

ninexnine_unit ninexnine_unit_3524(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W23000),
				.b1(W23010),
				.b2(W23020),
				.b3(W23100),
				.b4(W23110),
				.b5(W23120),
				.b6(W23200),
				.b7(W23210),
				.b8(W23220),
				.c(c20223)
);

ninexnine_unit ninexnine_unit_3525(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W23001),
				.b1(W23011),
				.b2(W23021),
				.b3(W23101),
				.b4(W23111),
				.b5(W23121),
				.b6(W23201),
				.b7(W23211),
				.b8(W23221),
				.c(c21223)
);

ninexnine_unit ninexnine_unit_3526(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W23002),
				.b1(W23012),
				.b2(W23022),
				.b3(W23102),
				.b4(W23112),
				.b5(W23122),
				.b6(W23202),
				.b7(W23212),
				.b8(W23222),
				.c(c22223)
);

ninexnine_unit ninexnine_unit_3527(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W23003),
				.b1(W23013),
				.b2(W23023),
				.b3(W23103),
				.b4(W23113),
				.b5(W23123),
				.b6(W23203),
				.b7(W23213),
				.b8(W23223),
				.c(c23223)
);

ninexnine_unit ninexnine_unit_3528(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W23004),
				.b1(W23014),
				.b2(W23024),
				.b3(W23104),
				.b4(W23114),
				.b5(W23124),
				.b6(W23204),
				.b7(W23214),
				.b8(W23224),
				.c(c24223)
);

ninexnine_unit ninexnine_unit_3529(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W23005),
				.b1(W23015),
				.b2(W23025),
				.b3(W23105),
				.b4(W23115),
				.b5(W23125),
				.b6(W23205),
				.b7(W23215),
				.b8(W23225),
				.c(c25223)
);

ninexnine_unit ninexnine_unit_3530(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W23006),
				.b1(W23016),
				.b2(W23026),
				.b3(W23106),
				.b4(W23116),
				.b5(W23126),
				.b6(W23206),
				.b7(W23216),
				.b8(W23226),
				.c(c26223)
);

ninexnine_unit ninexnine_unit_3531(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W23007),
				.b1(W23017),
				.b2(W23027),
				.b3(W23107),
				.b4(W23117),
				.b5(W23127),
				.b6(W23207),
				.b7(W23217),
				.b8(W23227),
				.c(c27223)
);

ninexnine_unit ninexnine_unit_3532(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W23008),
				.b1(W23018),
				.b2(W23028),
				.b3(W23108),
				.b4(W23118),
				.b5(W23128),
				.b6(W23208),
				.b7(W23218),
				.b8(W23228),
				.c(c28223)
);

ninexnine_unit ninexnine_unit_3533(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W23009),
				.b1(W23019),
				.b2(W23029),
				.b3(W23109),
				.b4(W23119),
				.b5(W23129),
				.b6(W23209),
				.b7(W23219),
				.b8(W23229),
				.c(c29223)
);

ninexnine_unit ninexnine_unit_3534(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2300A),
				.b1(W2301A),
				.b2(W2302A),
				.b3(W2310A),
				.b4(W2311A),
				.b5(W2312A),
				.b6(W2320A),
				.b7(W2321A),
				.b8(W2322A),
				.c(c2A223)
);

ninexnine_unit ninexnine_unit_3535(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2300B),
				.b1(W2301B),
				.b2(W2302B),
				.b3(W2310B),
				.b4(W2311B),
				.b5(W2312B),
				.b6(W2320B),
				.b7(W2321B),
				.b8(W2322B),
				.c(c2B223)
);

ninexnine_unit ninexnine_unit_3536(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2300C),
				.b1(W2301C),
				.b2(W2302C),
				.b3(W2310C),
				.b4(W2311C),
				.b5(W2312C),
				.b6(W2320C),
				.b7(W2321C),
				.b8(W2322C),
				.c(c2C223)
);

ninexnine_unit ninexnine_unit_3537(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2300D),
				.b1(W2301D),
				.b2(W2302D),
				.b3(W2310D),
				.b4(W2311D),
				.b5(W2312D),
				.b6(W2320D),
				.b7(W2321D),
				.b8(W2322D),
				.c(c2D223)
);

ninexnine_unit ninexnine_unit_3538(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2300E),
				.b1(W2301E),
				.b2(W2302E),
				.b3(W2310E),
				.b4(W2311E),
				.b5(W2312E),
				.b6(W2320E),
				.b7(W2321E),
				.b8(W2322E),
				.c(c2E223)
);

ninexnine_unit ninexnine_unit_3539(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2300F),
				.b1(W2301F),
				.b2(W2302F),
				.b3(W2310F),
				.b4(W2311F),
				.b5(W2312F),
				.b6(W2320F),
				.b7(W2321F),
				.b8(W2322F),
				.c(c2F223)
);

assign C2223=c20223+c21223+c22223+c23223+c24223+c25223+c26223+c27223+c28223+c29223+c2A223+c2B223+c2C223+c2D223+c2E223+c2F223;
assign A2223=(C2223>=0)?1:0;

assign P3223=A2223;

ninexnine_unit ninexnine_unit_3540(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20004)
);

ninexnine_unit ninexnine_unit_3541(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21004)
);

ninexnine_unit ninexnine_unit_3542(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22004)
);

ninexnine_unit ninexnine_unit_3543(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23004)
);

ninexnine_unit ninexnine_unit_3544(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24004)
);

ninexnine_unit ninexnine_unit_3545(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25004)
);

ninexnine_unit ninexnine_unit_3546(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26004)
);

ninexnine_unit ninexnine_unit_3547(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27004)
);

ninexnine_unit ninexnine_unit_3548(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W24008),
				.b1(W24018),
				.b2(W24028),
				.b3(W24108),
				.b4(W24118),
				.b5(W24128),
				.b6(W24208),
				.b7(W24218),
				.b8(W24228),
				.c(c28004)
);

ninexnine_unit ninexnine_unit_3549(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W24009),
				.b1(W24019),
				.b2(W24029),
				.b3(W24109),
				.b4(W24119),
				.b5(W24129),
				.b6(W24209),
				.b7(W24219),
				.b8(W24229),
				.c(c29004)
);

ninexnine_unit ninexnine_unit_3550(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2400A),
				.b1(W2401A),
				.b2(W2402A),
				.b3(W2410A),
				.b4(W2411A),
				.b5(W2412A),
				.b6(W2420A),
				.b7(W2421A),
				.b8(W2422A),
				.c(c2A004)
);

ninexnine_unit ninexnine_unit_3551(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2400B),
				.b1(W2401B),
				.b2(W2402B),
				.b3(W2410B),
				.b4(W2411B),
				.b5(W2412B),
				.b6(W2420B),
				.b7(W2421B),
				.b8(W2422B),
				.c(c2B004)
);

ninexnine_unit ninexnine_unit_3552(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2400C),
				.b1(W2401C),
				.b2(W2402C),
				.b3(W2410C),
				.b4(W2411C),
				.b5(W2412C),
				.b6(W2420C),
				.b7(W2421C),
				.b8(W2422C),
				.c(c2C004)
);

ninexnine_unit ninexnine_unit_3553(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2400D),
				.b1(W2401D),
				.b2(W2402D),
				.b3(W2410D),
				.b4(W2411D),
				.b5(W2412D),
				.b6(W2420D),
				.b7(W2421D),
				.b8(W2422D),
				.c(c2D004)
);

ninexnine_unit ninexnine_unit_3554(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2400E),
				.b1(W2401E),
				.b2(W2402E),
				.b3(W2410E),
				.b4(W2411E),
				.b5(W2412E),
				.b6(W2420E),
				.b7(W2421E),
				.b8(W2422E),
				.c(c2E004)
);

ninexnine_unit ninexnine_unit_3555(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2400F),
				.b1(W2401F),
				.b2(W2402F),
				.b3(W2410F),
				.b4(W2411F),
				.b5(W2412F),
				.b6(W2420F),
				.b7(W2421F),
				.b8(W2422F),
				.c(c2F004)
);

assign C2004=c20004+c21004+c22004+c23004+c24004+c25004+c26004+c27004+c28004+c29004+c2A004+c2B004+c2C004+c2D004+c2E004+c2F004;
assign A2004=(C2004>=0)?1:0;

assign P3004=A2004;

ninexnine_unit ninexnine_unit_3556(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20014)
);

ninexnine_unit ninexnine_unit_3557(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21014)
);

ninexnine_unit ninexnine_unit_3558(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22014)
);

ninexnine_unit ninexnine_unit_3559(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23014)
);

ninexnine_unit ninexnine_unit_3560(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24014)
);

ninexnine_unit ninexnine_unit_3561(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25014)
);

ninexnine_unit ninexnine_unit_3562(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26014)
);

ninexnine_unit ninexnine_unit_3563(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27014)
);

ninexnine_unit ninexnine_unit_3564(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W24008),
				.b1(W24018),
				.b2(W24028),
				.b3(W24108),
				.b4(W24118),
				.b5(W24128),
				.b6(W24208),
				.b7(W24218),
				.b8(W24228),
				.c(c28014)
);

ninexnine_unit ninexnine_unit_3565(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W24009),
				.b1(W24019),
				.b2(W24029),
				.b3(W24109),
				.b4(W24119),
				.b5(W24129),
				.b6(W24209),
				.b7(W24219),
				.b8(W24229),
				.c(c29014)
);

ninexnine_unit ninexnine_unit_3566(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2400A),
				.b1(W2401A),
				.b2(W2402A),
				.b3(W2410A),
				.b4(W2411A),
				.b5(W2412A),
				.b6(W2420A),
				.b7(W2421A),
				.b8(W2422A),
				.c(c2A014)
);

ninexnine_unit ninexnine_unit_3567(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2400B),
				.b1(W2401B),
				.b2(W2402B),
				.b3(W2410B),
				.b4(W2411B),
				.b5(W2412B),
				.b6(W2420B),
				.b7(W2421B),
				.b8(W2422B),
				.c(c2B014)
);

ninexnine_unit ninexnine_unit_3568(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2400C),
				.b1(W2401C),
				.b2(W2402C),
				.b3(W2410C),
				.b4(W2411C),
				.b5(W2412C),
				.b6(W2420C),
				.b7(W2421C),
				.b8(W2422C),
				.c(c2C014)
);

ninexnine_unit ninexnine_unit_3569(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2400D),
				.b1(W2401D),
				.b2(W2402D),
				.b3(W2410D),
				.b4(W2411D),
				.b5(W2412D),
				.b6(W2420D),
				.b7(W2421D),
				.b8(W2422D),
				.c(c2D014)
);

ninexnine_unit ninexnine_unit_3570(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2400E),
				.b1(W2401E),
				.b2(W2402E),
				.b3(W2410E),
				.b4(W2411E),
				.b5(W2412E),
				.b6(W2420E),
				.b7(W2421E),
				.b8(W2422E),
				.c(c2E014)
);

ninexnine_unit ninexnine_unit_3571(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2400F),
				.b1(W2401F),
				.b2(W2402F),
				.b3(W2410F),
				.b4(W2411F),
				.b5(W2412F),
				.b6(W2420F),
				.b7(W2421F),
				.b8(W2422F),
				.c(c2F014)
);

assign C2014=c20014+c21014+c22014+c23014+c24014+c25014+c26014+c27014+c28014+c29014+c2A014+c2B014+c2C014+c2D014+c2E014+c2F014;
assign A2014=(C2014>=0)?1:0;

assign P3014=A2014;

ninexnine_unit ninexnine_unit_3572(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20024)
);

ninexnine_unit ninexnine_unit_3573(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21024)
);

ninexnine_unit ninexnine_unit_3574(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22024)
);

ninexnine_unit ninexnine_unit_3575(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23024)
);

ninexnine_unit ninexnine_unit_3576(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24024)
);

ninexnine_unit ninexnine_unit_3577(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25024)
);

ninexnine_unit ninexnine_unit_3578(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26024)
);

ninexnine_unit ninexnine_unit_3579(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27024)
);

ninexnine_unit ninexnine_unit_3580(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W24008),
				.b1(W24018),
				.b2(W24028),
				.b3(W24108),
				.b4(W24118),
				.b5(W24128),
				.b6(W24208),
				.b7(W24218),
				.b8(W24228),
				.c(c28024)
);

ninexnine_unit ninexnine_unit_3581(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W24009),
				.b1(W24019),
				.b2(W24029),
				.b3(W24109),
				.b4(W24119),
				.b5(W24129),
				.b6(W24209),
				.b7(W24219),
				.b8(W24229),
				.c(c29024)
);

ninexnine_unit ninexnine_unit_3582(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2400A),
				.b1(W2401A),
				.b2(W2402A),
				.b3(W2410A),
				.b4(W2411A),
				.b5(W2412A),
				.b6(W2420A),
				.b7(W2421A),
				.b8(W2422A),
				.c(c2A024)
);

ninexnine_unit ninexnine_unit_3583(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2400B),
				.b1(W2401B),
				.b2(W2402B),
				.b3(W2410B),
				.b4(W2411B),
				.b5(W2412B),
				.b6(W2420B),
				.b7(W2421B),
				.b8(W2422B),
				.c(c2B024)
);

ninexnine_unit ninexnine_unit_3584(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2400C),
				.b1(W2401C),
				.b2(W2402C),
				.b3(W2410C),
				.b4(W2411C),
				.b5(W2412C),
				.b6(W2420C),
				.b7(W2421C),
				.b8(W2422C),
				.c(c2C024)
);

ninexnine_unit ninexnine_unit_3585(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2400D),
				.b1(W2401D),
				.b2(W2402D),
				.b3(W2410D),
				.b4(W2411D),
				.b5(W2412D),
				.b6(W2420D),
				.b7(W2421D),
				.b8(W2422D),
				.c(c2D024)
);

ninexnine_unit ninexnine_unit_3586(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2400E),
				.b1(W2401E),
				.b2(W2402E),
				.b3(W2410E),
				.b4(W2411E),
				.b5(W2412E),
				.b6(W2420E),
				.b7(W2421E),
				.b8(W2422E),
				.c(c2E024)
);

ninexnine_unit ninexnine_unit_3587(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2400F),
				.b1(W2401F),
				.b2(W2402F),
				.b3(W2410F),
				.b4(W2411F),
				.b5(W2412F),
				.b6(W2420F),
				.b7(W2421F),
				.b8(W2422F),
				.c(c2F024)
);

assign C2024=c20024+c21024+c22024+c23024+c24024+c25024+c26024+c27024+c28024+c29024+c2A024+c2B024+c2C024+c2D024+c2E024+c2F024;
assign A2024=(C2024>=0)?1:0;

assign P3024=A2024;

ninexnine_unit ninexnine_unit_3588(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20104)
);

ninexnine_unit ninexnine_unit_3589(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21104)
);

ninexnine_unit ninexnine_unit_3590(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22104)
);

ninexnine_unit ninexnine_unit_3591(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23104)
);

ninexnine_unit ninexnine_unit_3592(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24104)
);

ninexnine_unit ninexnine_unit_3593(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25104)
);

ninexnine_unit ninexnine_unit_3594(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26104)
);

ninexnine_unit ninexnine_unit_3595(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27104)
);

ninexnine_unit ninexnine_unit_3596(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W24008),
				.b1(W24018),
				.b2(W24028),
				.b3(W24108),
				.b4(W24118),
				.b5(W24128),
				.b6(W24208),
				.b7(W24218),
				.b8(W24228),
				.c(c28104)
);

ninexnine_unit ninexnine_unit_3597(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W24009),
				.b1(W24019),
				.b2(W24029),
				.b3(W24109),
				.b4(W24119),
				.b5(W24129),
				.b6(W24209),
				.b7(W24219),
				.b8(W24229),
				.c(c29104)
);

ninexnine_unit ninexnine_unit_3598(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2400A),
				.b1(W2401A),
				.b2(W2402A),
				.b3(W2410A),
				.b4(W2411A),
				.b5(W2412A),
				.b6(W2420A),
				.b7(W2421A),
				.b8(W2422A),
				.c(c2A104)
);

ninexnine_unit ninexnine_unit_3599(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2400B),
				.b1(W2401B),
				.b2(W2402B),
				.b3(W2410B),
				.b4(W2411B),
				.b5(W2412B),
				.b6(W2420B),
				.b7(W2421B),
				.b8(W2422B),
				.c(c2B104)
);

ninexnine_unit ninexnine_unit_3600(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2400C),
				.b1(W2401C),
				.b2(W2402C),
				.b3(W2410C),
				.b4(W2411C),
				.b5(W2412C),
				.b6(W2420C),
				.b7(W2421C),
				.b8(W2422C),
				.c(c2C104)
);

ninexnine_unit ninexnine_unit_3601(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2400D),
				.b1(W2401D),
				.b2(W2402D),
				.b3(W2410D),
				.b4(W2411D),
				.b5(W2412D),
				.b6(W2420D),
				.b7(W2421D),
				.b8(W2422D),
				.c(c2D104)
);

ninexnine_unit ninexnine_unit_3602(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2400E),
				.b1(W2401E),
				.b2(W2402E),
				.b3(W2410E),
				.b4(W2411E),
				.b5(W2412E),
				.b6(W2420E),
				.b7(W2421E),
				.b8(W2422E),
				.c(c2E104)
);

ninexnine_unit ninexnine_unit_3603(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2400F),
				.b1(W2401F),
				.b2(W2402F),
				.b3(W2410F),
				.b4(W2411F),
				.b5(W2412F),
				.b6(W2420F),
				.b7(W2421F),
				.b8(W2422F),
				.c(c2F104)
);

assign C2104=c20104+c21104+c22104+c23104+c24104+c25104+c26104+c27104+c28104+c29104+c2A104+c2B104+c2C104+c2D104+c2E104+c2F104;
assign A2104=(C2104>=0)?1:0;

assign P3104=A2104;

ninexnine_unit ninexnine_unit_3604(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20114)
);

ninexnine_unit ninexnine_unit_3605(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21114)
);

ninexnine_unit ninexnine_unit_3606(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22114)
);

ninexnine_unit ninexnine_unit_3607(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23114)
);

ninexnine_unit ninexnine_unit_3608(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24114)
);

ninexnine_unit ninexnine_unit_3609(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25114)
);

ninexnine_unit ninexnine_unit_3610(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26114)
);

ninexnine_unit ninexnine_unit_3611(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27114)
);

ninexnine_unit ninexnine_unit_3612(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W24008),
				.b1(W24018),
				.b2(W24028),
				.b3(W24108),
				.b4(W24118),
				.b5(W24128),
				.b6(W24208),
				.b7(W24218),
				.b8(W24228),
				.c(c28114)
);

ninexnine_unit ninexnine_unit_3613(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W24009),
				.b1(W24019),
				.b2(W24029),
				.b3(W24109),
				.b4(W24119),
				.b5(W24129),
				.b6(W24209),
				.b7(W24219),
				.b8(W24229),
				.c(c29114)
);

ninexnine_unit ninexnine_unit_3614(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2400A),
				.b1(W2401A),
				.b2(W2402A),
				.b3(W2410A),
				.b4(W2411A),
				.b5(W2412A),
				.b6(W2420A),
				.b7(W2421A),
				.b8(W2422A),
				.c(c2A114)
);

ninexnine_unit ninexnine_unit_3615(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2400B),
				.b1(W2401B),
				.b2(W2402B),
				.b3(W2410B),
				.b4(W2411B),
				.b5(W2412B),
				.b6(W2420B),
				.b7(W2421B),
				.b8(W2422B),
				.c(c2B114)
);

ninexnine_unit ninexnine_unit_3616(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2400C),
				.b1(W2401C),
				.b2(W2402C),
				.b3(W2410C),
				.b4(W2411C),
				.b5(W2412C),
				.b6(W2420C),
				.b7(W2421C),
				.b8(W2422C),
				.c(c2C114)
);

ninexnine_unit ninexnine_unit_3617(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2400D),
				.b1(W2401D),
				.b2(W2402D),
				.b3(W2410D),
				.b4(W2411D),
				.b5(W2412D),
				.b6(W2420D),
				.b7(W2421D),
				.b8(W2422D),
				.c(c2D114)
);

ninexnine_unit ninexnine_unit_3618(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2400E),
				.b1(W2401E),
				.b2(W2402E),
				.b3(W2410E),
				.b4(W2411E),
				.b5(W2412E),
				.b6(W2420E),
				.b7(W2421E),
				.b8(W2422E),
				.c(c2E114)
);

ninexnine_unit ninexnine_unit_3619(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2400F),
				.b1(W2401F),
				.b2(W2402F),
				.b3(W2410F),
				.b4(W2411F),
				.b5(W2412F),
				.b6(W2420F),
				.b7(W2421F),
				.b8(W2422F),
				.c(c2F114)
);

assign C2114=c20114+c21114+c22114+c23114+c24114+c25114+c26114+c27114+c28114+c29114+c2A114+c2B114+c2C114+c2D114+c2E114+c2F114;
assign A2114=(C2114>=0)?1:0;

assign P3114=A2114;

ninexnine_unit ninexnine_unit_3620(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20124)
);

ninexnine_unit ninexnine_unit_3621(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21124)
);

ninexnine_unit ninexnine_unit_3622(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22124)
);

ninexnine_unit ninexnine_unit_3623(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23124)
);

ninexnine_unit ninexnine_unit_3624(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24124)
);

ninexnine_unit ninexnine_unit_3625(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25124)
);

ninexnine_unit ninexnine_unit_3626(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26124)
);

ninexnine_unit ninexnine_unit_3627(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27124)
);

ninexnine_unit ninexnine_unit_3628(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W24008),
				.b1(W24018),
				.b2(W24028),
				.b3(W24108),
				.b4(W24118),
				.b5(W24128),
				.b6(W24208),
				.b7(W24218),
				.b8(W24228),
				.c(c28124)
);

ninexnine_unit ninexnine_unit_3629(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W24009),
				.b1(W24019),
				.b2(W24029),
				.b3(W24109),
				.b4(W24119),
				.b5(W24129),
				.b6(W24209),
				.b7(W24219),
				.b8(W24229),
				.c(c29124)
);

ninexnine_unit ninexnine_unit_3630(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2400A),
				.b1(W2401A),
				.b2(W2402A),
				.b3(W2410A),
				.b4(W2411A),
				.b5(W2412A),
				.b6(W2420A),
				.b7(W2421A),
				.b8(W2422A),
				.c(c2A124)
);

ninexnine_unit ninexnine_unit_3631(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2400B),
				.b1(W2401B),
				.b2(W2402B),
				.b3(W2410B),
				.b4(W2411B),
				.b5(W2412B),
				.b6(W2420B),
				.b7(W2421B),
				.b8(W2422B),
				.c(c2B124)
);

ninexnine_unit ninexnine_unit_3632(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2400C),
				.b1(W2401C),
				.b2(W2402C),
				.b3(W2410C),
				.b4(W2411C),
				.b5(W2412C),
				.b6(W2420C),
				.b7(W2421C),
				.b8(W2422C),
				.c(c2C124)
);

ninexnine_unit ninexnine_unit_3633(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2400D),
				.b1(W2401D),
				.b2(W2402D),
				.b3(W2410D),
				.b4(W2411D),
				.b5(W2412D),
				.b6(W2420D),
				.b7(W2421D),
				.b8(W2422D),
				.c(c2D124)
);

ninexnine_unit ninexnine_unit_3634(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2400E),
				.b1(W2401E),
				.b2(W2402E),
				.b3(W2410E),
				.b4(W2411E),
				.b5(W2412E),
				.b6(W2420E),
				.b7(W2421E),
				.b8(W2422E),
				.c(c2E124)
);

ninexnine_unit ninexnine_unit_3635(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2400F),
				.b1(W2401F),
				.b2(W2402F),
				.b3(W2410F),
				.b4(W2411F),
				.b5(W2412F),
				.b6(W2420F),
				.b7(W2421F),
				.b8(W2422F),
				.c(c2F124)
);

assign C2124=c20124+c21124+c22124+c23124+c24124+c25124+c26124+c27124+c28124+c29124+c2A124+c2B124+c2C124+c2D124+c2E124+c2F124;
assign A2124=(C2124>=0)?1:0;

assign P3124=A2124;

ninexnine_unit ninexnine_unit_3636(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20204)
);

ninexnine_unit ninexnine_unit_3637(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21204)
);

ninexnine_unit ninexnine_unit_3638(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22204)
);

ninexnine_unit ninexnine_unit_3639(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23204)
);

ninexnine_unit ninexnine_unit_3640(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24204)
);

ninexnine_unit ninexnine_unit_3641(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25204)
);

ninexnine_unit ninexnine_unit_3642(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26204)
);

ninexnine_unit ninexnine_unit_3643(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27204)
);

ninexnine_unit ninexnine_unit_3644(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W24008),
				.b1(W24018),
				.b2(W24028),
				.b3(W24108),
				.b4(W24118),
				.b5(W24128),
				.b6(W24208),
				.b7(W24218),
				.b8(W24228),
				.c(c28204)
);

ninexnine_unit ninexnine_unit_3645(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W24009),
				.b1(W24019),
				.b2(W24029),
				.b3(W24109),
				.b4(W24119),
				.b5(W24129),
				.b6(W24209),
				.b7(W24219),
				.b8(W24229),
				.c(c29204)
);

ninexnine_unit ninexnine_unit_3646(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2400A),
				.b1(W2401A),
				.b2(W2402A),
				.b3(W2410A),
				.b4(W2411A),
				.b5(W2412A),
				.b6(W2420A),
				.b7(W2421A),
				.b8(W2422A),
				.c(c2A204)
);

ninexnine_unit ninexnine_unit_3647(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2400B),
				.b1(W2401B),
				.b2(W2402B),
				.b3(W2410B),
				.b4(W2411B),
				.b5(W2412B),
				.b6(W2420B),
				.b7(W2421B),
				.b8(W2422B),
				.c(c2B204)
);

ninexnine_unit ninexnine_unit_3648(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2400C),
				.b1(W2401C),
				.b2(W2402C),
				.b3(W2410C),
				.b4(W2411C),
				.b5(W2412C),
				.b6(W2420C),
				.b7(W2421C),
				.b8(W2422C),
				.c(c2C204)
);

ninexnine_unit ninexnine_unit_3649(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2400D),
				.b1(W2401D),
				.b2(W2402D),
				.b3(W2410D),
				.b4(W2411D),
				.b5(W2412D),
				.b6(W2420D),
				.b7(W2421D),
				.b8(W2422D),
				.c(c2D204)
);

ninexnine_unit ninexnine_unit_3650(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2400E),
				.b1(W2401E),
				.b2(W2402E),
				.b3(W2410E),
				.b4(W2411E),
				.b5(W2412E),
				.b6(W2420E),
				.b7(W2421E),
				.b8(W2422E),
				.c(c2E204)
);

ninexnine_unit ninexnine_unit_3651(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2400F),
				.b1(W2401F),
				.b2(W2402F),
				.b3(W2410F),
				.b4(W2411F),
				.b5(W2412F),
				.b6(W2420F),
				.b7(W2421F),
				.b8(W2422F),
				.c(c2F204)
);

assign C2204=c20204+c21204+c22204+c23204+c24204+c25204+c26204+c27204+c28204+c29204+c2A204+c2B204+c2C204+c2D204+c2E204+c2F204;
assign A2204=(C2204>=0)?1:0;

assign P3204=A2204;

ninexnine_unit ninexnine_unit_3652(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20214)
);

ninexnine_unit ninexnine_unit_3653(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21214)
);

ninexnine_unit ninexnine_unit_3654(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22214)
);

ninexnine_unit ninexnine_unit_3655(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23214)
);

ninexnine_unit ninexnine_unit_3656(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24214)
);

ninexnine_unit ninexnine_unit_3657(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25214)
);

ninexnine_unit ninexnine_unit_3658(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26214)
);

ninexnine_unit ninexnine_unit_3659(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27214)
);

ninexnine_unit ninexnine_unit_3660(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W24008),
				.b1(W24018),
				.b2(W24028),
				.b3(W24108),
				.b4(W24118),
				.b5(W24128),
				.b6(W24208),
				.b7(W24218),
				.b8(W24228),
				.c(c28214)
);

ninexnine_unit ninexnine_unit_3661(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W24009),
				.b1(W24019),
				.b2(W24029),
				.b3(W24109),
				.b4(W24119),
				.b5(W24129),
				.b6(W24209),
				.b7(W24219),
				.b8(W24229),
				.c(c29214)
);

ninexnine_unit ninexnine_unit_3662(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2400A),
				.b1(W2401A),
				.b2(W2402A),
				.b3(W2410A),
				.b4(W2411A),
				.b5(W2412A),
				.b6(W2420A),
				.b7(W2421A),
				.b8(W2422A),
				.c(c2A214)
);

ninexnine_unit ninexnine_unit_3663(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2400B),
				.b1(W2401B),
				.b2(W2402B),
				.b3(W2410B),
				.b4(W2411B),
				.b5(W2412B),
				.b6(W2420B),
				.b7(W2421B),
				.b8(W2422B),
				.c(c2B214)
);

ninexnine_unit ninexnine_unit_3664(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2400C),
				.b1(W2401C),
				.b2(W2402C),
				.b3(W2410C),
				.b4(W2411C),
				.b5(W2412C),
				.b6(W2420C),
				.b7(W2421C),
				.b8(W2422C),
				.c(c2C214)
);

ninexnine_unit ninexnine_unit_3665(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2400D),
				.b1(W2401D),
				.b2(W2402D),
				.b3(W2410D),
				.b4(W2411D),
				.b5(W2412D),
				.b6(W2420D),
				.b7(W2421D),
				.b8(W2422D),
				.c(c2D214)
);

ninexnine_unit ninexnine_unit_3666(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2400E),
				.b1(W2401E),
				.b2(W2402E),
				.b3(W2410E),
				.b4(W2411E),
				.b5(W2412E),
				.b6(W2420E),
				.b7(W2421E),
				.b8(W2422E),
				.c(c2E214)
);

ninexnine_unit ninexnine_unit_3667(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2400F),
				.b1(W2401F),
				.b2(W2402F),
				.b3(W2410F),
				.b4(W2411F),
				.b5(W2412F),
				.b6(W2420F),
				.b7(W2421F),
				.b8(W2422F),
				.c(c2F214)
);

assign C2214=c20214+c21214+c22214+c23214+c24214+c25214+c26214+c27214+c28214+c29214+c2A214+c2B214+c2C214+c2D214+c2E214+c2F214;
assign A2214=(C2214>=0)?1:0;

assign P3214=A2214;

ninexnine_unit ninexnine_unit_3668(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W24000),
				.b1(W24010),
				.b2(W24020),
				.b3(W24100),
				.b4(W24110),
				.b5(W24120),
				.b6(W24200),
				.b7(W24210),
				.b8(W24220),
				.c(c20224)
);

ninexnine_unit ninexnine_unit_3669(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W24001),
				.b1(W24011),
				.b2(W24021),
				.b3(W24101),
				.b4(W24111),
				.b5(W24121),
				.b6(W24201),
				.b7(W24211),
				.b8(W24221),
				.c(c21224)
);

ninexnine_unit ninexnine_unit_3670(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W24002),
				.b1(W24012),
				.b2(W24022),
				.b3(W24102),
				.b4(W24112),
				.b5(W24122),
				.b6(W24202),
				.b7(W24212),
				.b8(W24222),
				.c(c22224)
);

ninexnine_unit ninexnine_unit_3671(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W24003),
				.b1(W24013),
				.b2(W24023),
				.b3(W24103),
				.b4(W24113),
				.b5(W24123),
				.b6(W24203),
				.b7(W24213),
				.b8(W24223),
				.c(c23224)
);

ninexnine_unit ninexnine_unit_3672(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W24004),
				.b1(W24014),
				.b2(W24024),
				.b3(W24104),
				.b4(W24114),
				.b5(W24124),
				.b6(W24204),
				.b7(W24214),
				.b8(W24224),
				.c(c24224)
);

ninexnine_unit ninexnine_unit_3673(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W24005),
				.b1(W24015),
				.b2(W24025),
				.b3(W24105),
				.b4(W24115),
				.b5(W24125),
				.b6(W24205),
				.b7(W24215),
				.b8(W24225),
				.c(c25224)
);

ninexnine_unit ninexnine_unit_3674(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W24006),
				.b1(W24016),
				.b2(W24026),
				.b3(W24106),
				.b4(W24116),
				.b5(W24126),
				.b6(W24206),
				.b7(W24216),
				.b8(W24226),
				.c(c26224)
);

ninexnine_unit ninexnine_unit_3675(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W24007),
				.b1(W24017),
				.b2(W24027),
				.b3(W24107),
				.b4(W24117),
				.b5(W24127),
				.b6(W24207),
				.b7(W24217),
				.b8(W24227),
				.c(c27224)
);

ninexnine_unit ninexnine_unit_3676(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W24008),
				.b1(W24018),
				.b2(W24028),
				.b3(W24108),
				.b4(W24118),
				.b5(W24128),
				.b6(W24208),
				.b7(W24218),
				.b8(W24228),
				.c(c28224)
);

ninexnine_unit ninexnine_unit_3677(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W24009),
				.b1(W24019),
				.b2(W24029),
				.b3(W24109),
				.b4(W24119),
				.b5(W24129),
				.b6(W24209),
				.b7(W24219),
				.b8(W24229),
				.c(c29224)
);

ninexnine_unit ninexnine_unit_3678(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2400A),
				.b1(W2401A),
				.b2(W2402A),
				.b3(W2410A),
				.b4(W2411A),
				.b5(W2412A),
				.b6(W2420A),
				.b7(W2421A),
				.b8(W2422A),
				.c(c2A224)
);

ninexnine_unit ninexnine_unit_3679(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2400B),
				.b1(W2401B),
				.b2(W2402B),
				.b3(W2410B),
				.b4(W2411B),
				.b5(W2412B),
				.b6(W2420B),
				.b7(W2421B),
				.b8(W2422B),
				.c(c2B224)
);

ninexnine_unit ninexnine_unit_3680(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2400C),
				.b1(W2401C),
				.b2(W2402C),
				.b3(W2410C),
				.b4(W2411C),
				.b5(W2412C),
				.b6(W2420C),
				.b7(W2421C),
				.b8(W2422C),
				.c(c2C224)
);

ninexnine_unit ninexnine_unit_3681(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2400D),
				.b1(W2401D),
				.b2(W2402D),
				.b3(W2410D),
				.b4(W2411D),
				.b5(W2412D),
				.b6(W2420D),
				.b7(W2421D),
				.b8(W2422D),
				.c(c2D224)
);

ninexnine_unit ninexnine_unit_3682(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2400E),
				.b1(W2401E),
				.b2(W2402E),
				.b3(W2410E),
				.b4(W2411E),
				.b5(W2412E),
				.b6(W2420E),
				.b7(W2421E),
				.b8(W2422E),
				.c(c2E224)
);

ninexnine_unit ninexnine_unit_3683(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2400F),
				.b1(W2401F),
				.b2(W2402F),
				.b3(W2410F),
				.b4(W2411F),
				.b5(W2412F),
				.b6(W2420F),
				.b7(W2421F),
				.b8(W2422F),
				.c(c2F224)
);

assign C2224=c20224+c21224+c22224+c23224+c24224+c25224+c26224+c27224+c28224+c29224+c2A224+c2B224+c2C224+c2D224+c2E224+c2F224;
assign A2224=(C2224>=0)?1:0;

assign P3224=A2224;

ninexnine_unit ninexnine_unit_3684(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20005)
);

ninexnine_unit ninexnine_unit_3685(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21005)
);

ninexnine_unit ninexnine_unit_3686(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22005)
);

ninexnine_unit ninexnine_unit_3687(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23005)
);

ninexnine_unit ninexnine_unit_3688(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24005)
);

ninexnine_unit ninexnine_unit_3689(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25005)
);

ninexnine_unit ninexnine_unit_3690(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26005)
);

ninexnine_unit ninexnine_unit_3691(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27005)
);

ninexnine_unit ninexnine_unit_3692(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W25008),
				.b1(W25018),
				.b2(W25028),
				.b3(W25108),
				.b4(W25118),
				.b5(W25128),
				.b6(W25208),
				.b7(W25218),
				.b8(W25228),
				.c(c28005)
);

ninexnine_unit ninexnine_unit_3693(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W25009),
				.b1(W25019),
				.b2(W25029),
				.b3(W25109),
				.b4(W25119),
				.b5(W25129),
				.b6(W25209),
				.b7(W25219),
				.b8(W25229),
				.c(c29005)
);

ninexnine_unit ninexnine_unit_3694(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2500A),
				.b1(W2501A),
				.b2(W2502A),
				.b3(W2510A),
				.b4(W2511A),
				.b5(W2512A),
				.b6(W2520A),
				.b7(W2521A),
				.b8(W2522A),
				.c(c2A005)
);

ninexnine_unit ninexnine_unit_3695(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2500B),
				.b1(W2501B),
				.b2(W2502B),
				.b3(W2510B),
				.b4(W2511B),
				.b5(W2512B),
				.b6(W2520B),
				.b7(W2521B),
				.b8(W2522B),
				.c(c2B005)
);

ninexnine_unit ninexnine_unit_3696(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2500C),
				.b1(W2501C),
				.b2(W2502C),
				.b3(W2510C),
				.b4(W2511C),
				.b5(W2512C),
				.b6(W2520C),
				.b7(W2521C),
				.b8(W2522C),
				.c(c2C005)
);

ninexnine_unit ninexnine_unit_3697(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2500D),
				.b1(W2501D),
				.b2(W2502D),
				.b3(W2510D),
				.b4(W2511D),
				.b5(W2512D),
				.b6(W2520D),
				.b7(W2521D),
				.b8(W2522D),
				.c(c2D005)
);

ninexnine_unit ninexnine_unit_3698(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2500E),
				.b1(W2501E),
				.b2(W2502E),
				.b3(W2510E),
				.b4(W2511E),
				.b5(W2512E),
				.b6(W2520E),
				.b7(W2521E),
				.b8(W2522E),
				.c(c2E005)
);

ninexnine_unit ninexnine_unit_3699(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2500F),
				.b1(W2501F),
				.b2(W2502F),
				.b3(W2510F),
				.b4(W2511F),
				.b5(W2512F),
				.b6(W2520F),
				.b7(W2521F),
				.b8(W2522F),
				.c(c2F005)
);

assign C2005=c20005+c21005+c22005+c23005+c24005+c25005+c26005+c27005+c28005+c29005+c2A005+c2B005+c2C005+c2D005+c2E005+c2F005;
assign A2005=(C2005>=0)?1:0;

assign P3005=A2005;

ninexnine_unit ninexnine_unit_3700(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20015)
);

ninexnine_unit ninexnine_unit_3701(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21015)
);

ninexnine_unit ninexnine_unit_3702(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22015)
);

ninexnine_unit ninexnine_unit_3703(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23015)
);

ninexnine_unit ninexnine_unit_3704(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24015)
);

ninexnine_unit ninexnine_unit_3705(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25015)
);

ninexnine_unit ninexnine_unit_3706(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26015)
);

ninexnine_unit ninexnine_unit_3707(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27015)
);

ninexnine_unit ninexnine_unit_3708(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W25008),
				.b1(W25018),
				.b2(W25028),
				.b3(W25108),
				.b4(W25118),
				.b5(W25128),
				.b6(W25208),
				.b7(W25218),
				.b8(W25228),
				.c(c28015)
);

ninexnine_unit ninexnine_unit_3709(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W25009),
				.b1(W25019),
				.b2(W25029),
				.b3(W25109),
				.b4(W25119),
				.b5(W25129),
				.b6(W25209),
				.b7(W25219),
				.b8(W25229),
				.c(c29015)
);

ninexnine_unit ninexnine_unit_3710(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2500A),
				.b1(W2501A),
				.b2(W2502A),
				.b3(W2510A),
				.b4(W2511A),
				.b5(W2512A),
				.b6(W2520A),
				.b7(W2521A),
				.b8(W2522A),
				.c(c2A015)
);

ninexnine_unit ninexnine_unit_3711(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2500B),
				.b1(W2501B),
				.b2(W2502B),
				.b3(W2510B),
				.b4(W2511B),
				.b5(W2512B),
				.b6(W2520B),
				.b7(W2521B),
				.b8(W2522B),
				.c(c2B015)
);

ninexnine_unit ninexnine_unit_3712(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2500C),
				.b1(W2501C),
				.b2(W2502C),
				.b3(W2510C),
				.b4(W2511C),
				.b5(W2512C),
				.b6(W2520C),
				.b7(W2521C),
				.b8(W2522C),
				.c(c2C015)
);

ninexnine_unit ninexnine_unit_3713(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2500D),
				.b1(W2501D),
				.b2(W2502D),
				.b3(W2510D),
				.b4(W2511D),
				.b5(W2512D),
				.b6(W2520D),
				.b7(W2521D),
				.b8(W2522D),
				.c(c2D015)
);

ninexnine_unit ninexnine_unit_3714(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2500E),
				.b1(W2501E),
				.b2(W2502E),
				.b3(W2510E),
				.b4(W2511E),
				.b5(W2512E),
				.b6(W2520E),
				.b7(W2521E),
				.b8(W2522E),
				.c(c2E015)
);

ninexnine_unit ninexnine_unit_3715(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2500F),
				.b1(W2501F),
				.b2(W2502F),
				.b3(W2510F),
				.b4(W2511F),
				.b5(W2512F),
				.b6(W2520F),
				.b7(W2521F),
				.b8(W2522F),
				.c(c2F015)
);

assign C2015=c20015+c21015+c22015+c23015+c24015+c25015+c26015+c27015+c28015+c29015+c2A015+c2B015+c2C015+c2D015+c2E015+c2F015;
assign A2015=(C2015>=0)?1:0;

assign P3015=A2015;

ninexnine_unit ninexnine_unit_3716(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20025)
);

ninexnine_unit ninexnine_unit_3717(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21025)
);

ninexnine_unit ninexnine_unit_3718(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22025)
);

ninexnine_unit ninexnine_unit_3719(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23025)
);

ninexnine_unit ninexnine_unit_3720(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24025)
);

ninexnine_unit ninexnine_unit_3721(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25025)
);

ninexnine_unit ninexnine_unit_3722(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26025)
);

ninexnine_unit ninexnine_unit_3723(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27025)
);

ninexnine_unit ninexnine_unit_3724(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W25008),
				.b1(W25018),
				.b2(W25028),
				.b3(W25108),
				.b4(W25118),
				.b5(W25128),
				.b6(W25208),
				.b7(W25218),
				.b8(W25228),
				.c(c28025)
);

ninexnine_unit ninexnine_unit_3725(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W25009),
				.b1(W25019),
				.b2(W25029),
				.b3(W25109),
				.b4(W25119),
				.b5(W25129),
				.b6(W25209),
				.b7(W25219),
				.b8(W25229),
				.c(c29025)
);

ninexnine_unit ninexnine_unit_3726(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2500A),
				.b1(W2501A),
				.b2(W2502A),
				.b3(W2510A),
				.b4(W2511A),
				.b5(W2512A),
				.b6(W2520A),
				.b7(W2521A),
				.b8(W2522A),
				.c(c2A025)
);

ninexnine_unit ninexnine_unit_3727(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2500B),
				.b1(W2501B),
				.b2(W2502B),
				.b3(W2510B),
				.b4(W2511B),
				.b5(W2512B),
				.b6(W2520B),
				.b7(W2521B),
				.b8(W2522B),
				.c(c2B025)
);

ninexnine_unit ninexnine_unit_3728(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2500C),
				.b1(W2501C),
				.b2(W2502C),
				.b3(W2510C),
				.b4(W2511C),
				.b5(W2512C),
				.b6(W2520C),
				.b7(W2521C),
				.b8(W2522C),
				.c(c2C025)
);

ninexnine_unit ninexnine_unit_3729(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2500D),
				.b1(W2501D),
				.b2(W2502D),
				.b3(W2510D),
				.b4(W2511D),
				.b5(W2512D),
				.b6(W2520D),
				.b7(W2521D),
				.b8(W2522D),
				.c(c2D025)
);

ninexnine_unit ninexnine_unit_3730(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2500E),
				.b1(W2501E),
				.b2(W2502E),
				.b3(W2510E),
				.b4(W2511E),
				.b5(W2512E),
				.b6(W2520E),
				.b7(W2521E),
				.b8(W2522E),
				.c(c2E025)
);

ninexnine_unit ninexnine_unit_3731(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2500F),
				.b1(W2501F),
				.b2(W2502F),
				.b3(W2510F),
				.b4(W2511F),
				.b5(W2512F),
				.b6(W2520F),
				.b7(W2521F),
				.b8(W2522F),
				.c(c2F025)
);

assign C2025=c20025+c21025+c22025+c23025+c24025+c25025+c26025+c27025+c28025+c29025+c2A025+c2B025+c2C025+c2D025+c2E025+c2F025;
assign A2025=(C2025>=0)?1:0;

assign P3025=A2025;

ninexnine_unit ninexnine_unit_3732(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20105)
);

ninexnine_unit ninexnine_unit_3733(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21105)
);

ninexnine_unit ninexnine_unit_3734(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22105)
);

ninexnine_unit ninexnine_unit_3735(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23105)
);

ninexnine_unit ninexnine_unit_3736(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24105)
);

ninexnine_unit ninexnine_unit_3737(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25105)
);

ninexnine_unit ninexnine_unit_3738(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26105)
);

ninexnine_unit ninexnine_unit_3739(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27105)
);

ninexnine_unit ninexnine_unit_3740(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W25008),
				.b1(W25018),
				.b2(W25028),
				.b3(W25108),
				.b4(W25118),
				.b5(W25128),
				.b6(W25208),
				.b7(W25218),
				.b8(W25228),
				.c(c28105)
);

ninexnine_unit ninexnine_unit_3741(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W25009),
				.b1(W25019),
				.b2(W25029),
				.b3(W25109),
				.b4(W25119),
				.b5(W25129),
				.b6(W25209),
				.b7(W25219),
				.b8(W25229),
				.c(c29105)
);

ninexnine_unit ninexnine_unit_3742(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2500A),
				.b1(W2501A),
				.b2(W2502A),
				.b3(W2510A),
				.b4(W2511A),
				.b5(W2512A),
				.b6(W2520A),
				.b7(W2521A),
				.b8(W2522A),
				.c(c2A105)
);

ninexnine_unit ninexnine_unit_3743(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2500B),
				.b1(W2501B),
				.b2(W2502B),
				.b3(W2510B),
				.b4(W2511B),
				.b5(W2512B),
				.b6(W2520B),
				.b7(W2521B),
				.b8(W2522B),
				.c(c2B105)
);

ninexnine_unit ninexnine_unit_3744(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2500C),
				.b1(W2501C),
				.b2(W2502C),
				.b3(W2510C),
				.b4(W2511C),
				.b5(W2512C),
				.b6(W2520C),
				.b7(W2521C),
				.b8(W2522C),
				.c(c2C105)
);

ninexnine_unit ninexnine_unit_3745(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2500D),
				.b1(W2501D),
				.b2(W2502D),
				.b3(W2510D),
				.b4(W2511D),
				.b5(W2512D),
				.b6(W2520D),
				.b7(W2521D),
				.b8(W2522D),
				.c(c2D105)
);

ninexnine_unit ninexnine_unit_3746(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2500E),
				.b1(W2501E),
				.b2(W2502E),
				.b3(W2510E),
				.b4(W2511E),
				.b5(W2512E),
				.b6(W2520E),
				.b7(W2521E),
				.b8(W2522E),
				.c(c2E105)
);

ninexnine_unit ninexnine_unit_3747(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2500F),
				.b1(W2501F),
				.b2(W2502F),
				.b3(W2510F),
				.b4(W2511F),
				.b5(W2512F),
				.b6(W2520F),
				.b7(W2521F),
				.b8(W2522F),
				.c(c2F105)
);

assign C2105=c20105+c21105+c22105+c23105+c24105+c25105+c26105+c27105+c28105+c29105+c2A105+c2B105+c2C105+c2D105+c2E105+c2F105;
assign A2105=(C2105>=0)?1:0;

assign P3105=A2105;

ninexnine_unit ninexnine_unit_3748(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20115)
);

ninexnine_unit ninexnine_unit_3749(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21115)
);

ninexnine_unit ninexnine_unit_3750(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22115)
);

ninexnine_unit ninexnine_unit_3751(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23115)
);

ninexnine_unit ninexnine_unit_3752(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24115)
);

ninexnine_unit ninexnine_unit_3753(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25115)
);

ninexnine_unit ninexnine_unit_3754(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26115)
);

ninexnine_unit ninexnine_unit_3755(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27115)
);

ninexnine_unit ninexnine_unit_3756(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W25008),
				.b1(W25018),
				.b2(W25028),
				.b3(W25108),
				.b4(W25118),
				.b5(W25128),
				.b6(W25208),
				.b7(W25218),
				.b8(W25228),
				.c(c28115)
);

ninexnine_unit ninexnine_unit_3757(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W25009),
				.b1(W25019),
				.b2(W25029),
				.b3(W25109),
				.b4(W25119),
				.b5(W25129),
				.b6(W25209),
				.b7(W25219),
				.b8(W25229),
				.c(c29115)
);

ninexnine_unit ninexnine_unit_3758(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2500A),
				.b1(W2501A),
				.b2(W2502A),
				.b3(W2510A),
				.b4(W2511A),
				.b5(W2512A),
				.b6(W2520A),
				.b7(W2521A),
				.b8(W2522A),
				.c(c2A115)
);

ninexnine_unit ninexnine_unit_3759(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2500B),
				.b1(W2501B),
				.b2(W2502B),
				.b3(W2510B),
				.b4(W2511B),
				.b5(W2512B),
				.b6(W2520B),
				.b7(W2521B),
				.b8(W2522B),
				.c(c2B115)
);

ninexnine_unit ninexnine_unit_3760(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2500C),
				.b1(W2501C),
				.b2(W2502C),
				.b3(W2510C),
				.b4(W2511C),
				.b5(W2512C),
				.b6(W2520C),
				.b7(W2521C),
				.b8(W2522C),
				.c(c2C115)
);

ninexnine_unit ninexnine_unit_3761(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2500D),
				.b1(W2501D),
				.b2(W2502D),
				.b3(W2510D),
				.b4(W2511D),
				.b5(W2512D),
				.b6(W2520D),
				.b7(W2521D),
				.b8(W2522D),
				.c(c2D115)
);

ninexnine_unit ninexnine_unit_3762(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2500E),
				.b1(W2501E),
				.b2(W2502E),
				.b3(W2510E),
				.b4(W2511E),
				.b5(W2512E),
				.b6(W2520E),
				.b7(W2521E),
				.b8(W2522E),
				.c(c2E115)
);

ninexnine_unit ninexnine_unit_3763(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2500F),
				.b1(W2501F),
				.b2(W2502F),
				.b3(W2510F),
				.b4(W2511F),
				.b5(W2512F),
				.b6(W2520F),
				.b7(W2521F),
				.b8(W2522F),
				.c(c2F115)
);

assign C2115=c20115+c21115+c22115+c23115+c24115+c25115+c26115+c27115+c28115+c29115+c2A115+c2B115+c2C115+c2D115+c2E115+c2F115;
assign A2115=(C2115>=0)?1:0;

assign P3115=A2115;

ninexnine_unit ninexnine_unit_3764(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20125)
);

ninexnine_unit ninexnine_unit_3765(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21125)
);

ninexnine_unit ninexnine_unit_3766(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22125)
);

ninexnine_unit ninexnine_unit_3767(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23125)
);

ninexnine_unit ninexnine_unit_3768(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24125)
);

ninexnine_unit ninexnine_unit_3769(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25125)
);

ninexnine_unit ninexnine_unit_3770(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26125)
);

ninexnine_unit ninexnine_unit_3771(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27125)
);

ninexnine_unit ninexnine_unit_3772(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W25008),
				.b1(W25018),
				.b2(W25028),
				.b3(W25108),
				.b4(W25118),
				.b5(W25128),
				.b6(W25208),
				.b7(W25218),
				.b8(W25228),
				.c(c28125)
);

ninexnine_unit ninexnine_unit_3773(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W25009),
				.b1(W25019),
				.b2(W25029),
				.b3(W25109),
				.b4(W25119),
				.b5(W25129),
				.b6(W25209),
				.b7(W25219),
				.b8(W25229),
				.c(c29125)
);

ninexnine_unit ninexnine_unit_3774(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2500A),
				.b1(W2501A),
				.b2(W2502A),
				.b3(W2510A),
				.b4(W2511A),
				.b5(W2512A),
				.b6(W2520A),
				.b7(W2521A),
				.b8(W2522A),
				.c(c2A125)
);

ninexnine_unit ninexnine_unit_3775(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2500B),
				.b1(W2501B),
				.b2(W2502B),
				.b3(W2510B),
				.b4(W2511B),
				.b5(W2512B),
				.b6(W2520B),
				.b7(W2521B),
				.b8(W2522B),
				.c(c2B125)
);

ninexnine_unit ninexnine_unit_3776(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2500C),
				.b1(W2501C),
				.b2(W2502C),
				.b3(W2510C),
				.b4(W2511C),
				.b5(W2512C),
				.b6(W2520C),
				.b7(W2521C),
				.b8(W2522C),
				.c(c2C125)
);

ninexnine_unit ninexnine_unit_3777(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2500D),
				.b1(W2501D),
				.b2(W2502D),
				.b3(W2510D),
				.b4(W2511D),
				.b5(W2512D),
				.b6(W2520D),
				.b7(W2521D),
				.b8(W2522D),
				.c(c2D125)
);

ninexnine_unit ninexnine_unit_3778(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2500E),
				.b1(W2501E),
				.b2(W2502E),
				.b3(W2510E),
				.b4(W2511E),
				.b5(W2512E),
				.b6(W2520E),
				.b7(W2521E),
				.b8(W2522E),
				.c(c2E125)
);

ninexnine_unit ninexnine_unit_3779(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2500F),
				.b1(W2501F),
				.b2(W2502F),
				.b3(W2510F),
				.b4(W2511F),
				.b5(W2512F),
				.b6(W2520F),
				.b7(W2521F),
				.b8(W2522F),
				.c(c2F125)
);

assign C2125=c20125+c21125+c22125+c23125+c24125+c25125+c26125+c27125+c28125+c29125+c2A125+c2B125+c2C125+c2D125+c2E125+c2F125;
assign A2125=(C2125>=0)?1:0;

assign P3125=A2125;

ninexnine_unit ninexnine_unit_3780(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20205)
);

ninexnine_unit ninexnine_unit_3781(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21205)
);

ninexnine_unit ninexnine_unit_3782(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22205)
);

ninexnine_unit ninexnine_unit_3783(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23205)
);

ninexnine_unit ninexnine_unit_3784(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24205)
);

ninexnine_unit ninexnine_unit_3785(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25205)
);

ninexnine_unit ninexnine_unit_3786(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26205)
);

ninexnine_unit ninexnine_unit_3787(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27205)
);

ninexnine_unit ninexnine_unit_3788(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W25008),
				.b1(W25018),
				.b2(W25028),
				.b3(W25108),
				.b4(W25118),
				.b5(W25128),
				.b6(W25208),
				.b7(W25218),
				.b8(W25228),
				.c(c28205)
);

ninexnine_unit ninexnine_unit_3789(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W25009),
				.b1(W25019),
				.b2(W25029),
				.b3(W25109),
				.b4(W25119),
				.b5(W25129),
				.b6(W25209),
				.b7(W25219),
				.b8(W25229),
				.c(c29205)
);

ninexnine_unit ninexnine_unit_3790(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2500A),
				.b1(W2501A),
				.b2(W2502A),
				.b3(W2510A),
				.b4(W2511A),
				.b5(W2512A),
				.b6(W2520A),
				.b7(W2521A),
				.b8(W2522A),
				.c(c2A205)
);

ninexnine_unit ninexnine_unit_3791(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2500B),
				.b1(W2501B),
				.b2(W2502B),
				.b3(W2510B),
				.b4(W2511B),
				.b5(W2512B),
				.b6(W2520B),
				.b7(W2521B),
				.b8(W2522B),
				.c(c2B205)
);

ninexnine_unit ninexnine_unit_3792(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2500C),
				.b1(W2501C),
				.b2(W2502C),
				.b3(W2510C),
				.b4(W2511C),
				.b5(W2512C),
				.b6(W2520C),
				.b7(W2521C),
				.b8(W2522C),
				.c(c2C205)
);

ninexnine_unit ninexnine_unit_3793(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2500D),
				.b1(W2501D),
				.b2(W2502D),
				.b3(W2510D),
				.b4(W2511D),
				.b5(W2512D),
				.b6(W2520D),
				.b7(W2521D),
				.b8(W2522D),
				.c(c2D205)
);

ninexnine_unit ninexnine_unit_3794(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2500E),
				.b1(W2501E),
				.b2(W2502E),
				.b3(W2510E),
				.b4(W2511E),
				.b5(W2512E),
				.b6(W2520E),
				.b7(W2521E),
				.b8(W2522E),
				.c(c2E205)
);

ninexnine_unit ninexnine_unit_3795(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2500F),
				.b1(W2501F),
				.b2(W2502F),
				.b3(W2510F),
				.b4(W2511F),
				.b5(W2512F),
				.b6(W2520F),
				.b7(W2521F),
				.b8(W2522F),
				.c(c2F205)
);

assign C2205=c20205+c21205+c22205+c23205+c24205+c25205+c26205+c27205+c28205+c29205+c2A205+c2B205+c2C205+c2D205+c2E205+c2F205;
assign A2205=(C2205>=0)?1:0;

assign P3205=A2205;

ninexnine_unit ninexnine_unit_3796(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20215)
);

ninexnine_unit ninexnine_unit_3797(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21215)
);

ninexnine_unit ninexnine_unit_3798(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22215)
);

ninexnine_unit ninexnine_unit_3799(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23215)
);

ninexnine_unit ninexnine_unit_3800(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24215)
);

ninexnine_unit ninexnine_unit_3801(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25215)
);

ninexnine_unit ninexnine_unit_3802(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26215)
);

ninexnine_unit ninexnine_unit_3803(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27215)
);

ninexnine_unit ninexnine_unit_3804(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W25008),
				.b1(W25018),
				.b2(W25028),
				.b3(W25108),
				.b4(W25118),
				.b5(W25128),
				.b6(W25208),
				.b7(W25218),
				.b8(W25228),
				.c(c28215)
);

ninexnine_unit ninexnine_unit_3805(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W25009),
				.b1(W25019),
				.b2(W25029),
				.b3(W25109),
				.b4(W25119),
				.b5(W25129),
				.b6(W25209),
				.b7(W25219),
				.b8(W25229),
				.c(c29215)
);

ninexnine_unit ninexnine_unit_3806(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2500A),
				.b1(W2501A),
				.b2(W2502A),
				.b3(W2510A),
				.b4(W2511A),
				.b5(W2512A),
				.b6(W2520A),
				.b7(W2521A),
				.b8(W2522A),
				.c(c2A215)
);

ninexnine_unit ninexnine_unit_3807(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2500B),
				.b1(W2501B),
				.b2(W2502B),
				.b3(W2510B),
				.b4(W2511B),
				.b5(W2512B),
				.b6(W2520B),
				.b7(W2521B),
				.b8(W2522B),
				.c(c2B215)
);

ninexnine_unit ninexnine_unit_3808(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2500C),
				.b1(W2501C),
				.b2(W2502C),
				.b3(W2510C),
				.b4(W2511C),
				.b5(W2512C),
				.b6(W2520C),
				.b7(W2521C),
				.b8(W2522C),
				.c(c2C215)
);

ninexnine_unit ninexnine_unit_3809(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2500D),
				.b1(W2501D),
				.b2(W2502D),
				.b3(W2510D),
				.b4(W2511D),
				.b5(W2512D),
				.b6(W2520D),
				.b7(W2521D),
				.b8(W2522D),
				.c(c2D215)
);

ninexnine_unit ninexnine_unit_3810(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2500E),
				.b1(W2501E),
				.b2(W2502E),
				.b3(W2510E),
				.b4(W2511E),
				.b5(W2512E),
				.b6(W2520E),
				.b7(W2521E),
				.b8(W2522E),
				.c(c2E215)
);

ninexnine_unit ninexnine_unit_3811(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2500F),
				.b1(W2501F),
				.b2(W2502F),
				.b3(W2510F),
				.b4(W2511F),
				.b5(W2512F),
				.b6(W2520F),
				.b7(W2521F),
				.b8(W2522F),
				.c(c2F215)
);

assign C2215=c20215+c21215+c22215+c23215+c24215+c25215+c26215+c27215+c28215+c29215+c2A215+c2B215+c2C215+c2D215+c2E215+c2F215;
assign A2215=(C2215>=0)?1:0;

assign P3215=A2215;

ninexnine_unit ninexnine_unit_3812(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W25000),
				.b1(W25010),
				.b2(W25020),
				.b3(W25100),
				.b4(W25110),
				.b5(W25120),
				.b6(W25200),
				.b7(W25210),
				.b8(W25220),
				.c(c20225)
);

ninexnine_unit ninexnine_unit_3813(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W25001),
				.b1(W25011),
				.b2(W25021),
				.b3(W25101),
				.b4(W25111),
				.b5(W25121),
				.b6(W25201),
				.b7(W25211),
				.b8(W25221),
				.c(c21225)
);

ninexnine_unit ninexnine_unit_3814(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W25002),
				.b1(W25012),
				.b2(W25022),
				.b3(W25102),
				.b4(W25112),
				.b5(W25122),
				.b6(W25202),
				.b7(W25212),
				.b8(W25222),
				.c(c22225)
);

ninexnine_unit ninexnine_unit_3815(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W25003),
				.b1(W25013),
				.b2(W25023),
				.b3(W25103),
				.b4(W25113),
				.b5(W25123),
				.b6(W25203),
				.b7(W25213),
				.b8(W25223),
				.c(c23225)
);

ninexnine_unit ninexnine_unit_3816(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W25004),
				.b1(W25014),
				.b2(W25024),
				.b3(W25104),
				.b4(W25114),
				.b5(W25124),
				.b6(W25204),
				.b7(W25214),
				.b8(W25224),
				.c(c24225)
);

ninexnine_unit ninexnine_unit_3817(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W25005),
				.b1(W25015),
				.b2(W25025),
				.b3(W25105),
				.b4(W25115),
				.b5(W25125),
				.b6(W25205),
				.b7(W25215),
				.b8(W25225),
				.c(c25225)
);

ninexnine_unit ninexnine_unit_3818(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W25006),
				.b1(W25016),
				.b2(W25026),
				.b3(W25106),
				.b4(W25116),
				.b5(W25126),
				.b6(W25206),
				.b7(W25216),
				.b8(W25226),
				.c(c26225)
);

ninexnine_unit ninexnine_unit_3819(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W25007),
				.b1(W25017),
				.b2(W25027),
				.b3(W25107),
				.b4(W25117),
				.b5(W25127),
				.b6(W25207),
				.b7(W25217),
				.b8(W25227),
				.c(c27225)
);

ninexnine_unit ninexnine_unit_3820(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W25008),
				.b1(W25018),
				.b2(W25028),
				.b3(W25108),
				.b4(W25118),
				.b5(W25128),
				.b6(W25208),
				.b7(W25218),
				.b8(W25228),
				.c(c28225)
);

ninexnine_unit ninexnine_unit_3821(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W25009),
				.b1(W25019),
				.b2(W25029),
				.b3(W25109),
				.b4(W25119),
				.b5(W25129),
				.b6(W25209),
				.b7(W25219),
				.b8(W25229),
				.c(c29225)
);

ninexnine_unit ninexnine_unit_3822(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2500A),
				.b1(W2501A),
				.b2(W2502A),
				.b3(W2510A),
				.b4(W2511A),
				.b5(W2512A),
				.b6(W2520A),
				.b7(W2521A),
				.b8(W2522A),
				.c(c2A225)
);

ninexnine_unit ninexnine_unit_3823(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2500B),
				.b1(W2501B),
				.b2(W2502B),
				.b3(W2510B),
				.b4(W2511B),
				.b5(W2512B),
				.b6(W2520B),
				.b7(W2521B),
				.b8(W2522B),
				.c(c2B225)
);

ninexnine_unit ninexnine_unit_3824(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2500C),
				.b1(W2501C),
				.b2(W2502C),
				.b3(W2510C),
				.b4(W2511C),
				.b5(W2512C),
				.b6(W2520C),
				.b7(W2521C),
				.b8(W2522C),
				.c(c2C225)
);

ninexnine_unit ninexnine_unit_3825(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2500D),
				.b1(W2501D),
				.b2(W2502D),
				.b3(W2510D),
				.b4(W2511D),
				.b5(W2512D),
				.b6(W2520D),
				.b7(W2521D),
				.b8(W2522D),
				.c(c2D225)
);

ninexnine_unit ninexnine_unit_3826(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2500E),
				.b1(W2501E),
				.b2(W2502E),
				.b3(W2510E),
				.b4(W2511E),
				.b5(W2512E),
				.b6(W2520E),
				.b7(W2521E),
				.b8(W2522E),
				.c(c2E225)
);

ninexnine_unit ninexnine_unit_3827(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2500F),
				.b1(W2501F),
				.b2(W2502F),
				.b3(W2510F),
				.b4(W2511F),
				.b5(W2512F),
				.b6(W2520F),
				.b7(W2521F),
				.b8(W2522F),
				.c(c2F225)
);

assign C2225=c20225+c21225+c22225+c23225+c24225+c25225+c26225+c27225+c28225+c29225+c2A225+c2B225+c2C225+c2D225+c2E225+c2F225;
assign A2225=(C2225>=0)?1:0;

assign P3225=A2225;

ninexnine_unit ninexnine_unit_3828(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20006)
);

ninexnine_unit ninexnine_unit_3829(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21006)
);

ninexnine_unit ninexnine_unit_3830(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22006)
);

ninexnine_unit ninexnine_unit_3831(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23006)
);

ninexnine_unit ninexnine_unit_3832(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24006)
);

ninexnine_unit ninexnine_unit_3833(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25006)
);

ninexnine_unit ninexnine_unit_3834(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26006)
);

ninexnine_unit ninexnine_unit_3835(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27006)
);

ninexnine_unit ninexnine_unit_3836(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W26008),
				.b1(W26018),
				.b2(W26028),
				.b3(W26108),
				.b4(W26118),
				.b5(W26128),
				.b6(W26208),
				.b7(W26218),
				.b8(W26228),
				.c(c28006)
);

ninexnine_unit ninexnine_unit_3837(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W26009),
				.b1(W26019),
				.b2(W26029),
				.b3(W26109),
				.b4(W26119),
				.b5(W26129),
				.b6(W26209),
				.b7(W26219),
				.b8(W26229),
				.c(c29006)
);

ninexnine_unit ninexnine_unit_3838(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2600A),
				.b1(W2601A),
				.b2(W2602A),
				.b3(W2610A),
				.b4(W2611A),
				.b5(W2612A),
				.b6(W2620A),
				.b7(W2621A),
				.b8(W2622A),
				.c(c2A006)
);

ninexnine_unit ninexnine_unit_3839(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2600B),
				.b1(W2601B),
				.b2(W2602B),
				.b3(W2610B),
				.b4(W2611B),
				.b5(W2612B),
				.b6(W2620B),
				.b7(W2621B),
				.b8(W2622B),
				.c(c2B006)
);

ninexnine_unit ninexnine_unit_3840(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2600C),
				.b1(W2601C),
				.b2(W2602C),
				.b3(W2610C),
				.b4(W2611C),
				.b5(W2612C),
				.b6(W2620C),
				.b7(W2621C),
				.b8(W2622C),
				.c(c2C006)
);

ninexnine_unit ninexnine_unit_3841(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2600D),
				.b1(W2601D),
				.b2(W2602D),
				.b3(W2610D),
				.b4(W2611D),
				.b5(W2612D),
				.b6(W2620D),
				.b7(W2621D),
				.b8(W2622D),
				.c(c2D006)
);

ninexnine_unit ninexnine_unit_3842(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2600E),
				.b1(W2601E),
				.b2(W2602E),
				.b3(W2610E),
				.b4(W2611E),
				.b5(W2612E),
				.b6(W2620E),
				.b7(W2621E),
				.b8(W2622E),
				.c(c2E006)
);

ninexnine_unit ninexnine_unit_3843(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2600F),
				.b1(W2601F),
				.b2(W2602F),
				.b3(W2610F),
				.b4(W2611F),
				.b5(W2612F),
				.b6(W2620F),
				.b7(W2621F),
				.b8(W2622F),
				.c(c2F006)
);

assign C2006=c20006+c21006+c22006+c23006+c24006+c25006+c26006+c27006+c28006+c29006+c2A006+c2B006+c2C006+c2D006+c2E006+c2F006;
assign A2006=(C2006>=0)?1:0;

assign P3006=A2006;

ninexnine_unit ninexnine_unit_3844(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20016)
);

ninexnine_unit ninexnine_unit_3845(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21016)
);

ninexnine_unit ninexnine_unit_3846(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22016)
);

ninexnine_unit ninexnine_unit_3847(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23016)
);

ninexnine_unit ninexnine_unit_3848(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24016)
);

ninexnine_unit ninexnine_unit_3849(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25016)
);

ninexnine_unit ninexnine_unit_3850(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26016)
);

ninexnine_unit ninexnine_unit_3851(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27016)
);

ninexnine_unit ninexnine_unit_3852(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W26008),
				.b1(W26018),
				.b2(W26028),
				.b3(W26108),
				.b4(W26118),
				.b5(W26128),
				.b6(W26208),
				.b7(W26218),
				.b8(W26228),
				.c(c28016)
);

ninexnine_unit ninexnine_unit_3853(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W26009),
				.b1(W26019),
				.b2(W26029),
				.b3(W26109),
				.b4(W26119),
				.b5(W26129),
				.b6(W26209),
				.b7(W26219),
				.b8(W26229),
				.c(c29016)
);

ninexnine_unit ninexnine_unit_3854(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2600A),
				.b1(W2601A),
				.b2(W2602A),
				.b3(W2610A),
				.b4(W2611A),
				.b5(W2612A),
				.b6(W2620A),
				.b7(W2621A),
				.b8(W2622A),
				.c(c2A016)
);

ninexnine_unit ninexnine_unit_3855(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2600B),
				.b1(W2601B),
				.b2(W2602B),
				.b3(W2610B),
				.b4(W2611B),
				.b5(W2612B),
				.b6(W2620B),
				.b7(W2621B),
				.b8(W2622B),
				.c(c2B016)
);

ninexnine_unit ninexnine_unit_3856(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2600C),
				.b1(W2601C),
				.b2(W2602C),
				.b3(W2610C),
				.b4(W2611C),
				.b5(W2612C),
				.b6(W2620C),
				.b7(W2621C),
				.b8(W2622C),
				.c(c2C016)
);

ninexnine_unit ninexnine_unit_3857(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2600D),
				.b1(W2601D),
				.b2(W2602D),
				.b3(W2610D),
				.b4(W2611D),
				.b5(W2612D),
				.b6(W2620D),
				.b7(W2621D),
				.b8(W2622D),
				.c(c2D016)
);

ninexnine_unit ninexnine_unit_3858(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2600E),
				.b1(W2601E),
				.b2(W2602E),
				.b3(W2610E),
				.b4(W2611E),
				.b5(W2612E),
				.b6(W2620E),
				.b7(W2621E),
				.b8(W2622E),
				.c(c2E016)
);

ninexnine_unit ninexnine_unit_3859(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2600F),
				.b1(W2601F),
				.b2(W2602F),
				.b3(W2610F),
				.b4(W2611F),
				.b5(W2612F),
				.b6(W2620F),
				.b7(W2621F),
				.b8(W2622F),
				.c(c2F016)
);

assign C2016=c20016+c21016+c22016+c23016+c24016+c25016+c26016+c27016+c28016+c29016+c2A016+c2B016+c2C016+c2D016+c2E016+c2F016;
assign A2016=(C2016>=0)?1:0;

assign P3016=A2016;

ninexnine_unit ninexnine_unit_3860(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20026)
);

ninexnine_unit ninexnine_unit_3861(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21026)
);

ninexnine_unit ninexnine_unit_3862(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22026)
);

ninexnine_unit ninexnine_unit_3863(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23026)
);

ninexnine_unit ninexnine_unit_3864(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24026)
);

ninexnine_unit ninexnine_unit_3865(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25026)
);

ninexnine_unit ninexnine_unit_3866(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26026)
);

ninexnine_unit ninexnine_unit_3867(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27026)
);

ninexnine_unit ninexnine_unit_3868(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W26008),
				.b1(W26018),
				.b2(W26028),
				.b3(W26108),
				.b4(W26118),
				.b5(W26128),
				.b6(W26208),
				.b7(W26218),
				.b8(W26228),
				.c(c28026)
);

ninexnine_unit ninexnine_unit_3869(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W26009),
				.b1(W26019),
				.b2(W26029),
				.b3(W26109),
				.b4(W26119),
				.b5(W26129),
				.b6(W26209),
				.b7(W26219),
				.b8(W26229),
				.c(c29026)
);

ninexnine_unit ninexnine_unit_3870(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2600A),
				.b1(W2601A),
				.b2(W2602A),
				.b3(W2610A),
				.b4(W2611A),
				.b5(W2612A),
				.b6(W2620A),
				.b7(W2621A),
				.b8(W2622A),
				.c(c2A026)
);

ninexnine_unit ninexnine_unit_3871(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2600B),
				.b1(W2601B),
				.b2(W2602B),
				.b3(W2610B),
				.b4(W2611B),
				.b5(W2612B),
				.b6(W2620B),
				.b7(W2621B),
				.b8(W2622B),
				.c(c2B026)
);

ninexnine_unit ninexnine_unit_3872(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2600C),
				.b1(W2601C),
				.b2(W2602C),
				.b3(W2610C),
				.b4(W2611C),
				.b5(W2612C),
				.b6(W2620C),
				.b7(W2621C),
				.b8(W2622C),
				.c(c2C026)
);

ninexnine_unit ninexnine_unit_3873(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2600D),
				.b1(W2601D),
				.b2(W2602D),
				.b3(W2610D),
				.b4(W2611D),
				.b5(W2612D),
				.b6(W2620D),
				.b7(W2621D),
				.b8(W2622D),
				.c(c2D026)
);

ninexnine_unit ninexnine_unit_3874(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2600E),
				.b1(W2601E),
				.b2(W2602E),
				.b3(W2610E),
				.b4(W2611E),
				.b5(W2612E),
				.b6(W2620E),
				.b7(W2621E),
				.b8(W2622E),
				.c(c2E026)
);

ninexnine_unit ninexnine_unit_3875(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2600F),
				.b1(W2601F),
				.b2(W2602F),
				.b3(W2610F),
				.b4(W2611F),
				.b5(W2612F),
				.b6(W2620F),
				.b7(W2621F),
				.b8(W2622F),
				.c(c2F026)
);

assign C2026=c20026+c21026+c22026+c23026+c24026+c25026+c26026+c27026+c28026+c29026+c2A026+c2B026+c2C026+c2D026+c2E026+c2F026;
assign A2026=(C2026>=0)?1:0;

assign P3026=A2026;

ninexnine_unit ninexnine_unit_3876(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20106)
);

ninexnine_unit ninexnine_unit_3877(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21106)
);

ninexnine_unit ninexnine_unit_3878(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22106)
);

ninexnine_unit ninexnine_unit_3879(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23106)
);

ninexnine_unit ninexnine_unit_3880(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24106)
);

ninexnine_unit ninexnine_unit_3881(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25106)
);

ninexnine_unit ninexnine_unit_3882(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26106)
);

ninexnine_unit ninexnine_unit_3883(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27106)
);

ninexnine_unit ninexnine_unit_3884(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W26008),
				.b1(W26018),
				.b2(W26028),
				.b3(W26108),
				.b4(W26118),
				.b5(W26128),
				.b6(W26208),
				.b7(W26218),
				.b8(W26228),
				.c(c28106)
);

ninexnine_unit ninexnine_unit_3885(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W26009),
				.b1(W26019),
				.b2(W26029),
				.b3(W26109),
				.b4(W26119),
				.b5(W26129),
				.b6(W26209),
				.b7(W26219),
				.b8(W26229),
				.c(c29106)
);

ninexnine_unit ninexnine_unit_3886(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2600A),
				.b1(W2601A),
				.b2(W2602A),
				.b3(W2610A),
				.b4(W2611A),
				.b5(W2612A),
				.b6(W2620A),
				.b7(W2621A),
				.b8(W2622A),
				.c(c2A106)
);

ninexnine_unit ninexnine_unit_3887(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2600B),
				.b1(W2601B),
				.b2(W2602B),
				.b3(W2610B),
				.b4(W2611B),
				.b5(W2612B),
				.b6(W2620B),
				.b7(W2621B),
				.b8(W2622B),
				.c(c2B106)
);

ninexnine_unit ninexnine_unit_3888(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2600C),
				.b1(W2601C),
				.b2(W2602C),
				.b3(W2610C),
				.b4(W2611C),
				.b5(W2612C),
				.b6(W2620C),
				.b7(W2621C),
				.b8(W2622C),
				.c(c2C106)
);

ninexnine_unit ninexnine_unit_3889(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2600D),
				.b1(W2601D),
				.b2(W2602D),
				.b3(W2610D),
				.b4(W2611D),
				.b5(W2612D),
				.b6(W2620D),
				.b7(W2621D),
				.b8(W2622D),
				.c(c2D106)
);

ninexnine_unit ninexnine_unit_3890(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2600E),
				.b1(W2601E),
				.b2(W2602E),
				.b3(W2610E),
				.b4(W2611E),
				.b5(W2612E),
				.b6(W2620E),
				.b7(W2621E),
				.b8(W2622E),
				.c(c2E106)
);

ninexnine_unit ninexnine_unit_3891(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2600F),
				.b1(W2601F),
				.b2(W2602F),
				.b3(W2610F),
				.b4(W2611F),
				.b5(W2612F),
				.b6(W2620F),
				.b7(W2621F),
				.b8(W2622F),
				.c(c2F106)
);

assign C2106=c20106+c21106+c22106+c23106+c24106+c25106+c26106+c27106+c28106+c29106+c2A106+c2B106+c2C106+c2D106+c2E106+c2F106;
assign A2106=(C2106>=0)?1:0;

assign P3106=A2106;

ninexnine_unit ninexnine_unit_3892(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20116)
);

ninexnine_unit ninexnine_unit_3893(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21116)
);

ninexnine_unit ninexnine_unit_3894(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22116)
);

ninexnine_unit ninexnine_unit_3895(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23116)
);

ninexnine_unit ninexnine_unit_3896(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24116)
);

ninexnine_unit ninexnine_unit_3897(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25116)
);

ninexnine_unit ninexnine_unit_3898(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26116)
);

ninexnine_unit ninexnine_unit_3899(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27116)
);

ninexnine_unit ninexnine_unit_3900(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W26008),
				.b1(W26018),
				.b2(W26028),
				.b3(W26108),
				.b4(W26118),
				.b5(W26128),
				.b6(W26208),
				.b7(W26218),
				.b8(W26228),
				.c(c28116)
);

ninexnine_unit ninexnine_unit_3901(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W26009),
				.b1(W26019),
				.b2(W26029),
				.b3(W26109),
				.b4(W26119),
				.b5(W26129),
				.b6(W26209),
				.b7(W26219),
				.b8(W26229),
				.c(c29116)
);

ninexnine_unit ninexnine_unit_3902(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2600A),
				.b1(W2601A),
				.b2(W2602A),
				.b3(W2610A),
				.b4(W2611A),
				.b5(W2612A),
				.b6(W2620A),
				.b7(W2621A),
				.b8(W2622A),
				.c(c2A116)
);

ninexnine_unit ninexnine_unit_3903(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2600B),
				.b1(W2601B),
				.b2(W2602B),
				.b3(W2610B),
				.b4(W2611B),
				.b5(W2612B),
				.b6(W2620B),
				.b7(W2621B),
				.b8(W2622B),
				.c(c2B116)
);

ninexnine_unit ninexnine_unit_3904(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2600C),
				.b1(W2601C),
				.b2(W2602C),
				.b3(W2610C),
				.b4(W2611C),
				.b5(W2612C),
				.b6(W2620C),
				.b7(W2621C),
				.b8(W2622C),
				.c(c2C116)
);

ninexnine_unit ninexnine_unit_3905(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2600D),
				.b1(W2601D),
				.b2(W2602D),
				.b3(W2610D),
				.b4(W2611D),
				.b5(W2612D),
				.b6(W2620D),
				.b7(W2621D),
				.b8(W2622D),
				.c(c2D116)
);

ninexnine_unit ninexnine_unit_3906(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2600E),
				.b1(W2601E),
				.b2(W2602E),
				.b3(W2610E),
				.b4(W2611E),
				.b5(W2612E),
				.b6(W2620E),
				.b7(W2621E),
				.b8(W2622E),
				.c(c2E116)
);

ninexnine_unit ninexnine_unit_3907(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2600F),
				.b1(W2601F),
				.b2(W2602F),
				.b3(W2610F),
				.b4(W2611F),
				.b5(W2612F),
				.b6(W2620F),
				.b7(W2621F),
				.b8(W2622F),
				.c(c2F116)
);

assign C2116=c20116+c21116+c22116+c23116+c24116+c25116+c26116+c27116+c28116+c29116+c2A116+c2B116+c2C116+c2D116+c2E116+c2F116;
assign A2116=(C2116>=0)?1:0;

assign P3116=A2116;

ninexnine_unit ninexnine_unit_3908(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20126)
);

ninexnine_unit ninexnine_unit_3909(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21126)
);

ninexnine_unit ninexnine_unit_3910(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22126)
);

ninexnine_unit ninexnine_unit_3911(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23126)
);

ninexnine_unit ninexnine_unit_3912(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24126)
);

ninexnine_unit ninexnine_unit_3913(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25126)
);

ninexnine_unit ninexnine_unit_3914(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26126)
);

ninexnine_unit ninexnine_unit_3915(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27126)
);

ninexnine_unit ninexnine_unit_3916(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W26008),
				.b1(W26018),
				.b2(W26028),
				.b3(W26108),
				.b4(W26118),
				.b5(W26128),
				.b6(W26208),
				.b7(W26218),
				.b8(W26228),
				.c(c28126)
);

ninexnine_unit ninexnine_unit_3917(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W26009),
				.b1(W26019),
				.b2(W26029),
				.b3(W26109),
				.b4(W26119),
				.b5(W26129),
				.b6(W26209),
				.b7(W26219),
				.b8(W26229),
				.c(c29126)
);

ninexnine_unit ninexnine_unit_3918(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2600A),
				.b1(W2601A),
				.b2(W2602A),
				.b3(W2610A),
				.b4(W2611A),
				.b5(W2612A),
				.b6(W2620A),
				.b7(W2621A),
				.b8(W2622A),
				.c(c2A126)
);

ninexnine_unit ninexnine_unit_3919(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2600B),
				.b1(W2601B),
				.b2(W2602B),
				.b3(W2610B),
				.b4(W2611B),
				.b5(W2612B),
				.b6(W2620B),
				.b7(W2621B),
				.b8(W2622B),
				.c(c2B126)
);

ninexnine_unit ninexnine_unit_3920(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2600C),
				.b1(W2601C),
				.b2(W2602C),
				.b3(W2610C),
				.b4(W2611C),
				.b5(W2612C),
				.b6(W2620C),
				.b7(W2621C),
				.b8(W2622C),
				.c(c2C126)
);

ninexnine_unit ninexnine_unit_3921(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2600D),
				.b1(W2601D),
				.b2(W2602D),
				.b3(W2610D),
				.b4(W2611D),
				.b5(W2612D),
				.b6(W2620D),
				.b7(W2621D),
				.b8(W2622D),
				.c(c2D126)
);

ninexnine_unit ninexnine_unit_3922(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2600E),
				.b1(W2601E),
				.b2(W2602E),
				.b3(W2610E),
				.b4(W2611E),
				.b5(W2612E),
				.b6(W2620E),
				.b7(W2621E),
				.b8(W2622E),
				.c(c2E126)
);

ninexnine_unit ninexnine_unit_3923(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2600F),
				.b1(W2601F),
				.b2(W2602F),
				.b3(W2610F),
				.b4(W2611F),
				.b5(W2612F),
				.b6(W2620F),
				.b7(W2621F),
				.b8(W2622F),
				.c(c2F126)
);

assign C2126=c20126+c21126+c22126+c23126+c24126+c25126+c26126+c27126+c28126+c29126+c2A126+c2B126+c2C126+c2D126+c2E126+c2F126;
assign A2126=(C2126>=0)?1:0;

assign P3126=A2126;

ninexnine_unit ninexnine_unit_3924(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20206)
);

ninexnine_unit ninexnine_unit_3925(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21206)
);

ninexnine_unit ninexnine_unit_3926(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22206)
);

ninexnine_unit ninexnine_unit_3927(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23206)
);

ninexnine_unit ninexnine_unit_3928(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24206)
);

ninexnine_unit ninexnine_unit_3929(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25206)
);

ninexnine_unit ninexnine_unit_3930(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26206)
);

ninexnine_unit ninexnine_unit_3931(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27206)
);

ninexnine_unit ninexnine_unit_3932(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W26008),
				.b1(W26018),
				.b2(W26028),
				.b3(W26108),
				.b4(W26118),
				.b5(W26128),
				.b6(W26208),
				.b7(W26218),
				.b8(W26228),
				.c(c28206)
);

ninexnine_unit ninexnine_unit_3933(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W26009),
				.b1(W26019),
				.b2(W26029),
				.b3(W26109),
				.b4(W26119),
				.b5(W26129),
				.b6(W26209),
				.b7(W26219),
				.b8(W26229),
				.c(c29206)
);

ninexnine_unit ninexnine_unit_3934(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2600A),
				.b1(W2601A),
				.b2(W2602A),
				.b3(W2610A),
				.b4(W2611A),
				.b5(W2612A),
				.b6(W2620A),
				.b7(W2621A),
				.b8(W2622A),
				.c(c2A206)
);

ninexnine_unit ninexnine_unit_3935(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2600B),
				.b1(W2601B),
				.b2(W2602B),
				.b3(W2610B),
				.b4(W2611B),
				.b5(W2612B),
				.b6(W2620B),
				.b7(W2621B),
				.b8(W2622B),
				.c(c2B206)
);

ninexnine_unit ninexnine_unit_3936(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2600C),
				.b1(W2601C),
				.b2(W2602C),
				.b3(W2610C),
				.b4(W2611C),
				.b5(W2612C),
				.b6(W2620C),
				.b7(W2621C),
				.b8(W2622C),
				.c(c2C206)
);

ninexnine_unit ninexnine_unit_3937(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2600D),
				.b1(W2601D),
				.b2(W2602D),
				.b3(W2610D),
				.b4(W2611D),
				.b5(W2612D),
				.b6(W2620D),
				.b7(W2621D),
				.b8(W2622D),
				.c(c2D206)
);

ninexnine_unit ninexnine_unit_3938(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2600E),
				.b1(W2601E),
				.b2(W2602E),
				.b3(W2610E),
				.b4(W2611E),
				.b5(W2612E),
				.b6(W2620E),
				.b7(W2621E),
				.b8(W2622E),
				.c(c2E206)
);

ninexnine_unit ninexnine_unit_3939(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2600F),
				.b1(W2601F),
				.b2(W2602F),
				.b3(W2610F),
				.b4(W2611F),
				.b5(W2612F),
				.b6(W2620F),
				.b7(W2621F),
				.b8(W2622F),
				.c(c2F206)
);

assign C2206=c20206+c21206+c22206+c23206+c24206+c25206+c26206+c27206+c28206+c29206+c2A206+c2B206+c2C206+c2D206+c2E206+c2F206;
assign A2206=(C2206>=0)?1:0;

assign P3206=A2206;

ninexnine_unit ninexnine_unit_3940(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20216)
);

ninexnine_unit ninexnine_unit_3941(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21216)
);

ninexnine_unit ninexnine_unit_3942(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22216)
);

ninexnine_unit ninexnine_unit_3943(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23216)
);

ninexnine_unit ninexnine_unit_3944(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24216)
);

ninexnine_unit ninexnine_unit_3945(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25216)
);

ninexnine_unit ninexnine_unit_3946(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26216)
);

ninexnine_unit ninexnine_unit_3947(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27216)
);

ninexnine_unit ninexnine_unit_3948(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W26008),
				.b1(W26018),
				.b2(W26028),
				.b3(W26108),
				.b4(W26118),
				.b5(W26128),
				.b6(W26208),
				.b7(W26218),
				.b8(W26228),
				.c(c28216)
);

ninexnine_unit ninexnine_unit_3949(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W26009),
				.b1(W26019),
				.b2(W26029),
				.b3(W26109),
				.b4(W26119),
				.b5(W26129),
				.b6(W26209),
				.b7(W26219),
				.b8(W26229),
				.c(c29216)
);

ninexnine_unit ninexnine_unit_3950(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2600A),
				.b1(W2601A),
				.b2(W2602A),
				.b3(W2610A),
				.b4(W2611A),
				.b5(W2612A),
				.b6(W2620A),
				.b7(W2621A),
				.b8(W2622A),
				.c(c2A216)
);

ninexnine_unit ninexnine_unit_3951(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2600B),
				.b1(W2601B),
				.b2(W2602B),
				.b3(W2610B),
				.b4(W2611B),
				.b5(W2612B),
				.b6(W2620B),
				.b7(W2621B),
				.b8(W2622B),
				.c(c2B216)
);

ninexnine_unit ninexnine_unit_3952(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2600C),
				.b1(W2601C),
				.b2(W2602C),
				.b3(W2610C),
				.b4(W2611C),
				.b5(W2612C),
				.b6(W2620C),
				.b7(W2621C),
				.b8(W2622C),
				.c(c2C216)
);

ninexnine_unit ninexnine_unit_3953(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2600D),
				.b1(W2601D),
				.b2(W2602D),
				.b3(W2610D),
				.b4(W2611D),
				.b5(W2612D),
				.b6(W2620D),
				.b7(W2621D),
				.b8(W2622D),
				.c(c2D216)
);

ninexnine_unit ninexnine_unit_3954(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2600E),
				.b1(W2601E),
				.b2(W2602E),
				.b3(W2610E),
				.b4(W2611E),
				.b5(W2612E),
				.b6(W2620E),
				.b7(W2621E),
				.b8(W2622E),
				.c(c2E216)
);

ninexnine_unit ninexnine_unit_3955(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2600F),
				.b1(W2601F),
				.b2(W2602F),
				.b3(W2610F),
				.b4(W2611F),
				.b5(W2612F),
				.b6(W2620F),
				.b7(W2621F),
				.b8(W2622F),
				.c(c2F216)
);

assign C2216=c20216+c21216+c22216+c23216+c24216+c25216+c26216+c27216+c28216+c29216+c2A216+c2B216+c2C216+c2D216+c2E216+c2F216;
assign A2216=(C2216>=0)?1:0;

assign P3216=A2216;

ninexnine_unit ninexnine_unit_3956(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W26000),
				.b1(W26010),
				.b2(W26020),
				.b3(W26100),
				.b4(W26110),
				.b5(W26120),
				.b6(W26200),
				.b7(W26210),
				.b8(W26220),
				.c(c20226)
);

ninexnine_unit ninexnine_unit_3957(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W26001),
				.b1(W26011),
				.b2(W26021),
				.b3(W26101),
				.b4(W26111),
				.b5(W26121),
				.b6(W26201),
				.b7(W26211),
				.b8(W26221),
				.c(c21226)
);

ninexnine_unit ninexnine_unit_3958(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W26002),
				.b1(W26012),
				.b2(W26022),
				.b3(W26102),
				.b4(W26112),
				.b5(W26122),
				.b6(W26202),
				.b7(W26212),
				.b8(W26222),
				.c(c22226)
);

ninexnine_unit ninexnine_unit_3959(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W26003),
				.b1(W26013),
				.b2(W26023),
				.b3(W26103),
				.b4(W26113),
				.b5(W26123),
				.b6(W26203),
				.b7(W26213),
				.b8(W26223),
				.c(c23226)
);

ninexnine_unit ninexnine_unit_3960(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W26004),
				.b1(W26014),
				.b2(W26024),
				.b3(W26104),
				.b4(W26114),
				.b5(W26124),
				.b6(W26204),
				.b7(W26214),
				.b8(W26224),
				.c(c24226)
);

ninexnine_unit ninexnine_unit_3961(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W26005),
				.b1(W26015),
				.b2(W26025),
				.b3(W26105),
				.b4(W26115),
				.b5(W26125),
				.b6(W26205),
				.b7(W26215),
				.b8(W26225),
				.c(c25226)
);

ninexnine_unit ninexnine_unit_3962(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W26006),
				.b1(W26016),
				.b2(W26026),
				.b3(W26106),
				.b4(W26116),
				.b5(W26126),
				.b6(W26206),
				.b7(W26216),
				.b8(W26226),
				.c(c26226)
);

ninexnine_unit ninexnine_unit_3963(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W26007),
				.b1(W26017),
				.b2(W26027),
				.b3(W26107),
				.b4(W26117),
				.b5(W26127),
				.b6(W26207),
				.b7(W26217),
				.b8(W26227),
				.c(c27226)
);

ninexnine_unit ninexnine_unit_3964(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W26008),
				.b1(W26018),
				.b2(W26028),
				.b3(W26108),
				.b4(W26118),
				.b5(W26128),
				.b6(W26208),
				.b7(W26218),
				.b8(W26228),
				.c(c28226)
);

ninexnine_unit ninexnine_unit_3965(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W26009),
				.b1(W26019),
				.b2(W26029),
				.b3(W26109),
				.b4(W26119),
				.b5(W26129),
				.b6(W26209),
				.b7(W26219),
				.b8(W26229),
				.c(c29226)
);

ninexnine_unit ninexnine_unit_3966(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2600A),
				.b1(W2601A),
				.b2(W2602A),
				.b3(W2610A),
				.b4(W2611A),
				.b5(W2612A),
				.b6(W2620A),
				.b7(W2621A),
				.b8(W2622A),
				.c(c2A226)
);

ninexnine_unit ninexnine_unit_3967(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2600B),
				.b1(W2601B),
				.b2(W2602B),
				.b3(W2610B),
				.b4(W2611B),
				.b5(W2612B),
				.b6(W2620B),
				.b7(W2621B),
				.b8(W2622B),
				.c(c2B226)
);

ninexnine_unit ninexnine_unit_3968(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2600C),
				.b1(W2601C),
				.b2(W2602C),
				.b3(W2610C),
				.b4(W2611C),
				.b5(W2612C),
				.b6(W2620C),
				.b7(W2621C),
				.b8(W2622C),
				.c(c2C226)
);

ninexnine_unit ninexnine_unit_3969(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2600D),
				.b1(W2601D),
				.b2(W2602D),
				.b3(W2610D),
				.b4(W2611D),
				.b5(W2612D),
				.b6(W2620D),
				.b7(W2621D),
				.b8(W2622D),
				.c(c2D226)
);

ninexnine_unit ninexnine_unit_3970(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2600E),
				.b1(W2601E),
				.b2(W2602E),
				.b3(W2610E),
				.b4(W2611E),
				.b5(W2612E),
				.b6(W2620E),
				.b7(W2621E),
				.b8(W2622E),
				.c(c2E226)
);

ninexnine_unit ninexnine_unit_3971(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2600F),
				.b1(W2601F),
				.b2(W2602F),
				.b3(W2610F),
				.b4(W2611F),
				.b5(W2612F),
				.b6(W2620F),
				.b7(W2621F),
				.b8(W2622F),
				.c(c2F226)
);

assign C2226=c20226+c21226+c22226+c23226+c24226+c25226+c26226+c27226+c28226+c29226+c2A226+c2B226+c2C226+c2D226+c2E226+c2F226;
assign A2226=(C2226>=0)?1:0;

assign P3226=A2226;

ninexnine_unit ninexnine_unit_3972(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20007)
);

ninexnine_unit ninexnine_unit_3973(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21007)
);

ninexnine_unit ninexnine_unit_3974(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22007)
);

ninexnine_unit ninexnine_unit_3975(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23007)
);

ninexnine_unit ninexnine_unit_3976(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24007)
);

ninexnine_unit ninexnine_unit_3977(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25007)
);

ninexnine_unit ninexnine_unit_3978(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26007)
);

ninexnine_unit ninexnine_unit_3979(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27007)
);

ninexnine_unit ninexnine_unit_3980(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W27008),
				.b1(W27018),
				.b2(W27028),
				.b3(W27108),
				.b4(W27118),
				.b5(W27128),
				.b6(W27208),
				.b7(W27218),
				.b8(W27228),
				.c(c28007)
);

ninexnine_unit ninexnine_unit_3981(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W27009),
				.b1(W27019),
				.b2(W27029),
				.b3(W27109),
				.b4(W27119),
				.b5(W27129),
				.b6(W27209),
				.b7(W27219),
				.b8(W27229),
				.c(c29007)
);

ninexnine_unit ninexnine_unit_3982(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2700A),
				.b1(W2701A),
				.b2(W2702A),
				.b3(W2710A),
				.b4(W2711A),
				.b5(W2712A),
				.b6(W2720A),
				.b7(W2721A),
				.b8(W2722A),
				.c(c2A007)
);

ninexnine_unit ninexnine_unit_3983(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2700B),
				.b1(W2701B),
				.b2(W2702B),
				.b3(W2710B),
				.b4(W2711B),
				.b5(W2712B),
				.b6(W2720B),
				.b7(W2721B),
				.b8(W2722B),
				.c(c2B007)
);

ninexnine_unit ninexnine_unit_3984(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2700C),
				.b1(W2701C),
				.b2(W2702C),
				.b3(W2710C),
				.b4(W2711C),
				.b5(W2712C),
				.b6(W2720C),
				.b7(W2721C),
				.b8(W2722C),
				.c(c2C007)
);

ninexnine_unit ninexnine_unit_3985(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2700D),
				.b1(W2701D),
				.b2(W2702D),
				.b3(W2710D),
				.b4(W2711D),
				.b5(W2712D),
				.b6(W2720D),
				.b7(W2721D),
				.b8(W2722D),
				.c(c2D007)
);

ninexnine_unit ninexnine_unit_3986(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2700E),
				.b1(W2701E),
				.b2(W2702E),
				.b3(W2710E),
				.b4(W2711E),
				.b5(W2712E),
				.b6(W2720E),
				.b7(W2721E),
				.b8(W2722E),
				.c(c2E007)
);

ninexnine_unit ninexnine_unit_3987(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2700F),
				.b1(W2701F),
				.b2(W2702F),
				.b3(W2710F),
				.b4(W2711F),
				.b5(W2712F),
				.b6(W2720F),
				.b7(W2721F),
				.b8(W2722F),
				.c(c2F007)
);

assign C2007=c20007+c21007+c22007+c23007+c24007+c25007+c26007+c27007+c28007+c29007+c2A007+c2B007+c2C007+c2D007+c2E007+c2F007;
assign A2007=(C2007>=0)?1:0;

assign P3007=A2007;

ninexnine_unit ninexnine_unit_3988(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20017)
);

ninexnine_unit ninexnine_unit_3989(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21017)
);

ninexnine_unit ninexnine_unit_3990(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22017)
);

ninexnine_unit ninexnine_unit_3991(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23017)
);

ninexnine_unit ninexnine_unit_3992(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24017)
);

ninexnine_unit ninexnine_unit_3993(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25017)
);

ninexnine_unit ninexnine_unit_3994(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26017)
);

ninexnine_unit ninexnine_unit_3995(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27017)
);

ninexnine_unit ninexnine_unit_3996(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W27008),
				.b1(W27018),
				.b2(W27028),
				.b3(W27108),
				.b4(W27118),
				.b5(W27128),
				.b6(W27208),
				.b7(W27218),
				.b8(W27228),
				.c(c28017)
);

ninexnine_unit ninexnine_unit_3997(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W27009),
				.b1(W27019),
				.b2(W27029),
				.b3(W27109),
				.b4(W27119),
				.b5(W27129),
				.b6(W27209),
				.b7(W27219),
				.b8(W27229),
				.c(c29017)
);

ninexnine_unit ninexnine_unit_3998(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2700A),
				.b1(W2701A),
				.b2(W2702A),
				.b3(W2710A),
				.b4(W2711A),
				.b5(W2712A),
				.b6(W2720A),
				.b7(W2721A),
				.b8(W2722A),
				.c(c2A017)
);

ninexnine_unit ninexnine_unit_3999(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2700B),
				.b1(W2701B),
				.b2(W2702B),
				.b3(W2710B),
				.b4(W2711B),
				.b5(W2712B),
				.b6(W2720B),
				.b7(W2721B),
				.b8(W2722B),
				.c(c2B017)
);

ninexnine_unit ninexnine_unit_4000(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2700C),
				.b1(W2701C),
				.b2(W2702C),
				.b3(W2710C),
				.b4(W2711C),
				.b5(W2712C),
				.b6(W2720C),
				.b7(W2721C),
				.b8(W2722C),
				.c(c2C017)
);

ninexnine_unit ninexnine_unit_4001(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2700D),
				.b1(W2701D),
				.b2(W2702D),
				.b3(W2710D),
				.b4(W2711D),
				.b5(W2712D),
				.b6(W2720D),
				.b7(W2721D),
				.b8(W2722D),
				.c(c2D017)
);

ninexnine_unit ninexnine_unit_4002(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2700E),
				.b1(W2701E),
				.b2(W2702E),
				.b3(W2710E),
				.b4(W2711E),
				.b5(W2712E),
				.b6(W2720E),
				.b7(W2721E),
				.b8(W2722E),
				.c(c2E017)
);

ninexnine_unit ninexnine_unit_4003(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2700F),
				.b1(W2701F),
				.b2(W2702F),
				.b3(W2710F),
				.b4(W2711F),
				.b5(W2712F),
				.b6(W2720F),
				.b7(W2721F),
				.b8(W2722F),
				.c(c2F017)
);

assign C2017=c20017+c21017+c22017+c23017+c24017+c25017+c26017+c27017+c28017+c29017+c2A017+c2B017+c2C017+c2D017+c2E017+c2F017;
assign A2017=(C2017>=0)?1:0;

assign P3017=A2017;

ninexnine_unit ninexnine_unit_4004(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20027)
);

ninexnine_unit ninexnine_unit_4005(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21027)
);

ninexnine_unit ninexnine_unit_4006(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22027)
);

ninexnine_unit ninexnine_unit_4007(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23027)
);

ninexnine_unit ninexnine_unit_4008(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24027)
);

ninexnine_unit ninexnine_unit_4009(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25027)
);

ninexnine_unit ninexnine_unit_4010(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26027)
);

ninexnine_unit ninexnine_unit_4011(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27027)
);

ninexnine_unit ninexnine_unit_4012(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W27008),
				.b1(W27018),
				.b2(W27028),
				.b3(W27108),
				.b4(W27118),
				.b5(W27128),
				.b6(W27208),
				.b7(W27218),
				.b8(W27228),
				.c(c28027)
);

ninexnine_unit ninexnine_unit_4013(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W27009),
				.b1(W27019),
				.b2(W27029),
				.b3(W27109),
				.b4(W27119),
				.b5(W27129),
				.b6(W27209),
				.b7(W27219),
				.b8(W27229),
				.c(c29027)
);

ninexnine_unit ninexnine_unit_4014(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2700A),
				.b1(W2701A),
				.b2(W2702A),
				.b3(W2710A),
				.b4(W2711A),
				.b5(W2712A),
				.b6(W2720A),
				.b7(W2721A),
				.b8(W2722A),
				.c(c2A027)
);

ninexnine_unit ninexnine_unit_4015(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2700B),
				.b1(W2701B),
				.b2(W2702B),
				.b3(W2710B),
				.b4(W2711B),
				.b5(W2712B),
				.b6(W2720B),
				.b7(W2721B),
				.b8(W2722B),
				.c(c2B027)
);

ninexnine_unit ninexnine_unit_4016(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2700C),
				.b1(W2701C),
				.b2(W2702C),
				.b3(W2710C),
				.b4(W2711C),
				.b5(W2712C),
				.b6(W2720C),
				.b7(W2721C),
				.b8(W2722C),
				.c(c2C027)
);

ninexnine_unit ninexnine_unit_4017(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2700D),
				.b1(W2701D),
				.b2(W2702D),
				.b3(W2710D),
				.b4(W2711D),
				.b5(W2712D),
				.b6(W2720D),
				.b7(W2721D),
				.b8(W2722D),
				.c(c2D027)
);

ninexnine_unit ninexnine_unit_4018(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2700E),
				.b1(W2701E),
				.b2(W2702E),
				.b3(W2710E),
				.b4(W2711E),
				.b5(W2712E),
				.b6(W2720E),
				.b7(W2721E),
				.b8(W2722E),
				.c(c2E027)
);

ninexnine_unit ninexnine_unit_4019(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2700F),
				.b1(W2701F),
				.b2(W2702F),
				.b3(W2710F),
				.b4(W2711F),
				.b5(W2712F),
				.b6(W2720F),
				.b7(W2721F),
				.b8(W2722F),
				.c(c2F027)
);

assign C2027=c20027+c21027+c22027+c23027+c24027+c25027+c26027+c27027+c28027+c29027+c2A027+c2B027+c2C027+c2D027+c2E027+c2F027;
assign A2027=(C2027>=0)?1:0;

assign P3027=A2027;

ninexnine_unit ninexnine_unit_4020(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20107)
);

ninexnine_unit ninexnine_unit_4021(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21107)
);

ninexnine_unit ninexnine_unit_4022(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22107)
);

ninexnine_unit ninexnine_unit_4023(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23107)
);

ninexnine_unit ninexnine_unit_4024(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24107)
);

ninexnine_unit ninexnine_unit_4025(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25107)
);

ninexnine_unit ninexnine_unit_4026(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26107)
);

ninexnine_unit ninexnine_unit_4027(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27107)
);

ninexnine_unit ninexnine_unit_4028(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W27008),
				.b1(W27018),
				.b2(W27028),
				.b3(W27108),
				.b4(W27118),
				.b5(W27128),
				.b6(W27208),
				.b7(W27218),
				.b8(W27228),
				.c(c28107)
);

ninexnine_unit ninexnine_unit_4029(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W27009),
				.b1(W27019),
				.b2(W27029),
				.b3(W27109),
				.b4(W27119),
				.b5(W27129),
				.b6(W27209),
				.b7(W27219),
				.b8(W27229),
				.c(c29107)
);

ninexnine_unit ninexnine_unit_4030(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2700A),
				.b1(W2701A),
				.b2(W2702A),
				.b3(W2710A),
				.b4(W2711A),
				.b5(W2712A),
				.b6(W2720A),
				.b7(W2721A),
				.b8(W2722A),
				.c(c2A107)
);

ninexnine_unit ninexnine_unit_4031(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2700B),
				.b1(W2701B),
				.b2(W2702B),
				.b3(W2710B),
				.b4(W2711B),
				.b5(W2712B),
				.b6(W2720B),
				.b7(W2721B),
				.b8(W2722B),
				.c(c2B107)
);

ninexnine_unit ninexnine_unit_4032(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2700C),
				.b1(W2701C),
				.b2(W2702C),
				.b3(W2710C),
				.b4(W2711C),
				.b5(W2712C),
				.b6(W2720C),
				.b7(W2721C),
				.b8(W2722C),
				.c(c2C107)
);

ninexnine_unit ninexnine_unit_4033(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2700D),
				.b1(W2701D),
				.b2(W2702D),
				.b3(W2710D),
				.b4(W2711D),
				.b5(W2712D),
				.b6(W2720D),
				.b7(W2721D),
				.b8(W2722D),
				.c(c2D107)
);

ninexnine_unit ninexnine_unit_4034(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2700E),
				.b1(W2701E),
				.b2(W2702E),
				.b3(W2710E),
				.b4(W2711E),
				.b5(W2712E),
				.b6(W2720E),
				.b7(W2721E),
				.b8(W2722E),
				.c(c2E107)
);

ninexnine_unit ninexnine_unit_4035(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2700F),
				.b1(W2701F),
				.b2(W2702F),
				.b3(W2710F),
				.b4(W2711F),
				.b5(W2712F),
				.b6(W2720F),
				.b7(W2721F),
				.b8(W2722F),
				.c(c2F107)
);

assign C2107=c20107+c21107+c22107+c23107+c24107+c25107+c26107+c27107+c28107+c29107+c2A107+c2B107+c2C107+c2D107+c2E107+c2F107;
assign A2107=(C2107>=0)?1:0;

assign P3107=A2107;

ninexnine_unit ninexnine_unit_4036(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20117)
);

ninexnine_unit ninexnine_unit_4037(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21117)
);

ninexnine_unit ninexnine_unit_4038(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22117)
);

ninexnine_unit ninexnine_unit_4039(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23117)
);

ninexnine_unit ninexnine_unit_4040(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24117)
);

ninexnine_unit ninexnine_unit_4041(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25117)
);

ninexnine_unit ninexnine_unit_4042(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26117)
);

ninexnine_unit ninexnine_unit_4043(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27117)
);

ninexnine_unit ninexnine_unit_4044(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W27008),
				.b1(W27018),
				.b2(W27028),
				.b3(W27108),
				.b4(W27118),
				.b5(W27128),
				.b6(W27208),
				.b7(W27218),
				.b8(W27228),
				.c(c28117)
);

ninexnine_unit ninexnine_unit_4045(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W27009),
				.b1(W27019),
				.b2(W27029),
				.b3(W27109),
				.b4(W27119),
				.b5(W27129),
				.b6(W27209),
				.b7(W27219),
				.b8(W27229),
				.c(c29117)
);

ninexnine_unit ninexnine_unit_4046(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2700A),
				.b1(W2701A),
				.b2(W2702A),
				.b3(W2710A),
				.b4(W2711A),
				.b5(W2712A),
				.b6(W2720A),
				.b7(W2721A),
				.b8(W2722A),
				.c(c2A117)
);

ninexnine_unit ninexnine_unit_4047(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2700B),
				.b1(W2701B),
				.b2(W2702B),
				.b3(W2710B),
				.b4(W2711B),
				.b5(W2712B),
				.b6(W2720B),
				.b7(W2721B),
				.b8(W2722B),
				.c(c2B117)
);

ninexnine_unit ninexnine_unit_4048(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2700C),
				.b1(W2701C),
				.b2(W2702C),
				.b3(W2710C),
				.b4(W2711C),
				.b5(W2712C),
				.b6(W2720C),
				.b7(W2721C),
				.b8(W2722C),
				.c(c2C117)
);

ninexnine_unit ninexnine_unit_4049(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2700D),
				.b1(W2701D),
				.b2(W2702D),
				.b3(W2710D),
				.b4(W2711D),
				.b5(W2712D),
				.b6(W2720D),
				.b7(W2721D),
				.b8(W2722D),
				.c(c2D117)
);

ninexnine_unit ninexnine_unit_4050(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2700E),
				.b1(W2701E),
				.b2(W2702E),
				.b3(W2710E),
				.b4(W2711E),
				.b5(W2712E),
				.b6(W2720E),
				.b7(W2721E),
				.b8(W2722E),
				.c(c2E117)
);

ninexnine_unit ninexnine_unit_4051(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2700F),
				.b1(W2701F),
				.b2(W2702F),
				.b3(W2710F),
				.b4(W2711F),
				.b5(W2712F),
				.b6(W2720F),
				.b7(W2721F),
				.b8(W2722F),
				.c(c2F117)
);

assign C2117=c20117+c21117+c22117+c23117+c24117+c25117+c26117+c27117+c28117+c29117+c2A117+c2B117+c2C117+c2D117+c2E117+c2F117;
assign A2117=(C2117>=0)?1:0;

assign P3117=A2117;

ninexnine_unit ninexnine_unit_4052(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20127)
);

ninexnine_unit ninexnine_unit_4053(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21127)
);

ninexnine_unit ninexnine_unit_4054(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22127)
);

ninexnine_unit ninexnine_unit_4055(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23127)
);

ninexnine_unit ninexnine_unit_4056(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24127)
);

ninexnine_unit ninexnine_unit_4057(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25127)
);

ninexnine_unit ninexnine_unit_4058(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26127)
);

ninexnine_unit ninexnine_unit_4059(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27127)
);

ninexnine_unit ninexnine_unit_4060(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W27008),
				.b1(W27018),
				.b2(W27028),
				.b3(W27108),
				.b4(W27118),
				.b5(W27128),
				.b6(W27208),
				.b7(W27218),
				.b8(W27228),
				.c(c28127)
);

ninexnine_unit ninexnine_unit_4061(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W27009),
				.b1(W27019),
				.b2(W27029),
				.b3(W27109),
				.b4(W27119),
				.b5(W27129),
				.b6(W27209),
				.b7(W27219),
				.b8(W27229),
				.c(c29127)
);

ninexnine_unit ninexnine_unit_4062(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2700A),
				.b1(W2701A),
				.b2(W2702A),
				.b3(W2710A),
				.b4(W2711A),
				.b5(W2712A),
				.b6(W2720A),
				.b7(W2721A),
				.b8(W2722A),
				.c(c2A127)
);

ninexnine_unit ninexnine_unit_4063(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2700B),
				.b1(W2701B),
				.b2(W2702B),
				.b3(W2710B),
				.b4(W2711B),
				.b5(W2712B),
				.b6(W2720B),
				.b7(W2721B),
				.b8(W2722B),
				.c(c2B127)
);

ninexnine_unit ninexnine_unit_4064(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2700C),
				.b1(W2701C),
				.b2(W2702C),
				.b3(W2710C),
				.b4(W2711C),
				.b5(W2712C),
				.b6(W2720C),
				.b7(W2721C),
				.b8(W2722C),
				.c(c2C127)
);

ninexnine_unit ninexnine_unit_4065(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2700D),
				.b1(W2701D),
				.b2(W2702D),
				.b3(W2710D),
				.b4(W2711D),
				.b5(W2712D),
				.b6(W2720D),
				.b7(W2721D),
				.b8(W2722D),
				.c(c2D127)
);

ninexnine_unit ninexnine_unit_4066(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2700E),
				.b1(W2701E),
				.b2(W2702E),
				.b3(W2710E),
				.b4(W2711E),
				.b5(W2712E),
				.b6(W2720E),
				.b7(W2721E),
				.b8(W2722E),
				.c(c2E127)
);

ninexnine_unit ninexnine_unit_4067(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2700F),
				.b1(W2701F),
				.b2(W2702F),
				.b3(W2710F),
				.b4(W2711F),
				.b5(W2712F),
				.b6(W2720F),
				.b7(W2721F),
				.b8(W2722F),
				.c(c2F127)
);

assign C2127=c20127+c21127+c22127+c23127+c24127+c25127+c26127+c27127+c28127+c29127+c2A127+c2B127+c2C127+c2D127+c2E127+c2F127;
assign A2127=(C2127>=0)?1:0;

assign P3127=A2127;

ninexnine_unit ninexnine_unit_4068(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20207)
);

ninexnine_unit ninexnine_unit_4069(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21207)
);

ninexnine_unit ninexnine_unit_4070(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22207)
);

ninexnine_unit ninexnine_unit_4071(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23207)
);

ninexnine_unit ninexnine_unit_4072(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24207)
);

ninexnine_unit ninexnine_unit_4073(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25207)
);

ninexnine_unit ninexnine_unit_4074(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26207)
);

ninexnine_unit ninexnine_unit_4075(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27207)
);

ninexnine_unit ninexnine_unit_4076(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W27008),
				.b1(W27018),
				.b2(W27028),
				.b3(W27108),
				.b4(W27118),
				.b5(W27128),
				.b6(W27208),
				.b7(W27218),
				.b8(W27228),
				.c(c28207)
);

ninexnine_unit ninexnine_unit_4077(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W27009),
				.b1(W27019),
				.b2(W27029),
				.b3(W27109),
				.b4(W27119),
				.b5(W27129),
				.b6(W27209),
				.b7(W27219),
				.b8(W27229),
				.c(c29207)
);

ninexnine_unit ninexnine_unit_4078(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2700A),
				.b1(W2701A),
				.b2(W2702A),
				.b3(W2710A),
				.b4(W2711A),
				.b5(W2712A),
				.b6(W2720A),
				.b7(W2721A),
				.b8(W2722A),
				.c(c2A207)
);

ninexnine_unit ninexnine_unit_4079(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2700B),
				.b1(W2701B),
				.b2(W2702B),
				.b3(W2710B),
				.b4(W2711B),
				.b5(W2712B),
				.b6(W2720B),
				.b7(W2721B),
				.b8(W2722B),
				.c(c2B207)
);

ninexnine_unit ninexnine_unit_4080(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2700C),
				.b1(W2701C),
				.b2(W2702C),
				.b3(W2710C),
				.b4(W2711C),
				.b5(W2712C),
				.b6(W2720C),
				.b7(W2721C),
				.b8(W2722C),
				.c(c2C207)
);

ninexnine_unit ninexnine_unit_4081(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2700D),
				.b1(W2701D),
				.b2(W2702D),
				.b3(W2710D),
				.b4(W2711D),
				.b5(W2712D),
				.b6(W2720D),
				.b7(W2721D),
				.b8(W2722D),
				.c(c2D207)
);

ninexnine_unit ninexnine_unit_4082(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2700E),
				.b1(W2701E),
				.b2(W2702E),
				.b3(W2710E),
				.b4(W2711E),
				.b5(W2712E),
				.b6(W2720E),
				.b7(W2721E),
				.b8(W2722E),
				.c(c2E207)
);

ninexnine_unit ninexnine_unit_4083(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2700F),
				.b1(W2701F),
				.b2(W2702F),
				.b3(W2710F),
				.b4(W2711F),
				.b5(W2712F),
				.b6(W2720F),
				.b7(W2721F),
				.b8(W2722F),
				.c(c2F207)
);

assign C2207=c20207+c21207+c22207+c23207+c24207+c25207+c26207+c27207+c28207+c29207+c2A207+c2B207+c2C207+c2D207+c2E207+c2F207;
assign A2207=(C2207>=0)?1:0;

assign P3207=A2207;

ninexnine_unit ninexnine_unit_4084(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20217)
);

ninexnine_unit ninexnine_unit_4085(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21217)
);

ninexnine_unit ninexnine_unit_4086(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22217)
);

ninexnine_unit ninexnine_unit_4087(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23217)
);

ninexnine_unit ninexnine_unit_4088(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24217)
);

ninexnine_unit ninexnine_unit_4089(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25217)
);

ninexnine_unit ninexnine_unit_4090(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26217)
);

ninexnine_unit ninexnine_unit_4091(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27217)
);

ninexnine_unit ninexnine_unit_4092(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W27008),
				.b1(W27018),
				.b2(W27028),
				.b3(W27108),
				.b4(W27118),
				.b5(W27128),
				.b6(W27208),
				.b7(W27218),
				.b8(W27228),
				.c(c28217)
);

ninexnine_unit ninexnine_unit_4093(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W27009),
				.b1(W27019),
				.b2(W27029),
				.b3(W27109),
				.b4(W27119),
				.b5(W27129),
				.b6(W27209),
				.b7(W27219),
				.b8(W27229),
				.c(c29217)
);

ninexnine_unit ninexnine_unit_4094(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2700A),
				.b1(W2701A),
				.b2(W2702A),
				.b3(W2710A),
				.b4(W2711A),
				.b5(W2712A),
				.b6(W2720A),
				.b7(W2721A),
				.b8(W2722A),
				.c(c2A217)
);

ninexnine_unit ninexnine_unit_4095(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2700B),
				.b1(W2701B),
				.b2(W2702B),
				.b3(W2710B),
				.b4(W2711B),
				.b5(W2712B),
				.b6(W2720B),
				.b7(W2721B),
				.b8(W2722B),
				.c(c2B217)
);

ninexnine_unit ninexnine_unit_4096(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2700C),
				.b1(W2701C),
				.b2(W2702C),
				.b3(W2710C),
				.b4(W2711C),
				.b5(W2712C),
				.b6(W2720C),
				.b7(W2721C),
				.b8(W2722C),
				.c(c2C217)
);

ninexnine_unit ninexnine_unit_4097(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2700D),
				.b1(W2701D),
				.b2(W2702D),
				.b3(W2710D),
				.b4(W2711D),
				.b5(W2712D),
				.b6(W2720D),
				.b7(W2721D),
				.b8(W2722D),
				.c(c2D217)
);

ninexnine_unit ninexnine_unit_4098(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2700E),
				.b1(W2701E),
				.b2(W2702E),
				.b3(W2710E),
				.b4(W2711E),
				.b5(W2712E),
				.b6(W2720E),
				.b7(W2721E),
				.b8(W2722E),
				.c(c2E217)
);

ninexnine_unit ninexnine_unit_4099(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2700F),
				.b1(W2701F),
				.b2(W2702F),
				.b3(W2710F),
				.b4(W2711F),
				.b5(W2712F),
				.b6(W2720F),
				.b7(W2721F),
				.b8(W2722F),
				.c(c2F217)
);

assign C2217=c20217+c21217+c22217+c23217+c24217+c25217+c26217+c27217+c28217+c29217+c2A217+c2B217+c2C217+c2D217+c2E217+c2F217;
assign A2217=(C2217>=0)?1:0;

assign P3217=A2217;

ninexnine_unit ninexnine_unit_4100(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W27000),
				.b1(W27010),
				.b2(W27020),
				.b3(W27100),
				.b4(W27110),
				.b5(W27120),
				.b6(W27200),
				.b7(W27210),
				.b8(W27220),
				.c(c20227)
);

ninexnine_unit ninexnine_unit_4101(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W27001),
				.b1(W27011),
				.b2(W27021),
				.b3(W27101),
				.b4(W27111),
				.b5(W27121),
				.b6(W27201),
				.b7(W27211),
				.b8(W27221),
				.c(c21227)
);

ninexnine_unit ninexnine_unit_4102(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W27002),
				.b1(W27012),
				.b2(W27022),
				.b3(W27102),
				.b4(W27112),
				.b5(W27122),
				.b6(W27202),
				.b7(W27212),
				.b8(W27222),
				.c(c22227)
);

ninexnine_unit ninexnine_unit_4103(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W27003),
				.b1(W27013),
				.b2(W27023),
				.b3(W27103),
				.b4(W27113),
				.b5(W27123),
				.b6(W27203),
				.b7(W27213),
				.b8(W27223),
				.c(c23227)
);

ninexnine_unit ninexnine_unit_4104(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W27004),
				.b1(W27014),
				.b2(W27024),
				.b3(W27104),
				.b4(W27114),
				.b5(W27124),
				.b6(W27204),
				.b7(W27214),
				.b8(W27224),
				.c(c24227)
);

ninexnine_unit ninexnine_unit_4105(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W27005),
				.b1(W27015),
				.b2(W27025),
				.b3(W27105),
				.b4(W27115),
				.b5(W27125),
				.b6(W27205),
				.b7(W27215),
				.b8(W27225),
				.c(c25227)
);

ninexnine_unit ninexnine_unit_4106(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W27006),
				.b1(W27016),
				.b2(W27026),
				.b3(W27106),
				.b4(W27116),
				.b5(W27126),
				.b6(W27206),
				.b7(W27216),
				.b8(W27226),
				.c(c26227)
);

ninexnine_unit ninexnine_unit_4107(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W27007),
				.b1(W27017),
				.b2(W27027),
				.b3(W27107),
				.b4(W27117),
				.b5(W27127),
				.b6(W27207),
				.b7(W27217),
				.b8(W27227),
				.c(c27227)
);

ninexnine_unit ninexnine_unit_4108(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W27008),
				.b1(W27018),
				.b2(W27028),
				.b3(W27108),
				.b4(W27118),
				.b5(W27128),
				.b6(W27208),
				.b7(W27218),
				.b8(W27228),
				.c(c28227)
);

ninexnine_unit ninexnine_unit_4109(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W27009),
				.b1(W27019),
				.b2(W27029),
				.b3(W27109),
				.b4(W27119),
				.b5(W27129),
				.b6(W27209),
				.b7(W27219),
				.b8(W27229),
				.c(c29227)
);

ninexnine_unit ninexnine_unit_4110(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2700A),
				.b1(W2701A),
				.b2(W2702A),
				.b3(W2710A),
				.b4(W2711A),
				.b5(W2712A),
				.b6(W2720A),
				.b7(W2721A),
				.b8(W2722A),
				.c(c2A227)
);

ninexnine_unit ninexnine_unit_4111(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2700B),
				.b1(W2701B),
				.b2(W2702B),
				.b3(W2710B),
				.b4(W2711B),
				.b5(W2712B),
				.b6(W2720B),
				.b7(W2721B),
				.b8(W2722B),
				.c(c2B227)
);

ninexnine_unit ninexnine_unit_4112(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2700C),
				.b1(W2701C),
				.b2(W2702C),
				.b3(W2710C),
				.b4(W2711C),
				.b5(W2712C),
				.b6(W2720C),
				.b7(W2721C),
				.b8(W2722C),
				.c(c2C227)
);

ninexnine_unit ninexnine_unit_4113(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2700D),
				.b1(W2701D),
				.b2(W2702D),
				.b3(W2710D),
				.b4(W2711D),
				.b5(W2712D),
				.b6(W2720D),
				.b7(W2721D),
				.b8(W2722D),
				.c(c2D227)
);

ninexnine_unit ninexnine_unit_4114(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2700E),
				.b1(W2701E),
				.b2(W2702E),
				.b3(W2710E),
				.b4(W2711E),
				.b5(W2712E),
				.b6(W2720E),
				.b7(W2721E),
				.b8(W2722E),
				.c(c2E227)
);

ninexnine_unit ninexnine_unit_4115(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2700F),
				.b1(W2701F),
				.b2(W2702F),
				.b3(W2710F),
				.b4(W2711F),
				.b5(W2712F),
				.b6(W2720F),
				.b7(W2721F),
				.b8(W2722F),
				.c(c2F227)
);

assign C2227=c20227+c21227+c22227+c23227+c24227+c25227+c26227+c27227+c28227+c29227+c2A227+c2B227+c2C227+c2D227+c2E227+c2F227;
assign A2227=(C2227>=0)?1:0;

assign P3227=A2227;

ninexnine_unit ninexnine_unit_4116(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20008)
);

ninexnine_unit ninexnine_unit_4117(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21008)
);

ninexnine_unit ninexnine_unit_4118(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22008)
);

ninexnine_unit ninexnine_unit_4119(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23008)
);

ninexnine_unit ninexnine_unit_4120(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24008)
);

ninexnine_unit ninexnine_unit_4121(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25008)
);

ninexnine_unit ninexnine_unit_4122(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26008)
);

ninexnine_unit ninexnine_unit_4123(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27008)
);

ninexnine_unit ninexnine_unit_4124(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W28008),
				.b1(W28018),
				.b2(W28028),
				.b3(W28108),
				.b4(W28118),
				.b5(W28128),
				.b6(W28208),
				.b7(W28218),
				.b8(W28228),
				.c(c28008)
);

ninexnine_unit ninexnine_unit_4125(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W28009),
				.b1(W28019),
				.b2(W28029),
				.b3(W28109),
				.b4(W28119),
				.b5(W28129),
				.b6(W28209),
				.b7(W28219),
				.b8(W28229),
				.c(c29008)
);

ninexnine_unit ninexnine_unit_4126(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2800A),
				.b1(W2801A),
				.b2(W2802A),
				.b3(W2810A),
				.b4(W2811A),
				.b5(W2812A),
				.b6(W2820A),
				.b7(W2821A),
				.b8(W2822A),
				.c(c2A008)
);

ninexnine_unit ninexnine_unit_4127(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2800B),
				.b1(W2801B),
				.b2(W2802B),
				.b3(W2810B),
				.b4(W2811B),
				.b5(W2812B),
				.b6(W2820B),
				.b7(W2821B),
				.b8(W2822B),
				.c(c2B008)
);

ninexnine_unit ninexnine_unit_4128(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2800C),
				.b1(W2801C),
				.b2(W2802C),
				.b3(W2810C),
				.b4(W2811C),
				.b5(W2812C),
				.b6(W2820C),
				.b7(W2821C),
				.b8(W2822C),
				.c(c2C008)
);

ninexnine_unit ninexnine_unit_4129(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2800D),
				.b1(W2801D),
				.b2(W2802D),
				.b3(W2810D),
				.b4(W2811D),
				.b5(W2812D),
				.b6(W2820D),
				.b7(W2821D),
				.b8(W2822D),
				.c(c2D008)
);

ninexnine_unit ninexnine_unit_4130(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2800E),
				.b1(W2801E),
				.b2(W2802E),
				.b3(W2810E),
				.b4(W2811E),
				.b5(W2812E),
				.b6(W2820E),
				.b7(W2821E),
				.b8(W2822E),
				.c(c2E008)
);

ninexnine_unit ninexnine_unit_4131(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2800F),
				.b1(W2801F),
				.b2(W2802F),
				.b3(W2810F),
				.b4(W2811F),
				.b5(W2812F),
				.b6(W2820F),
				.b7(W2821F),
				.b8(W2822F),
				.c(c2F008)
);

assign C2008=c20008+c21008+c22008+c23008+c24008+c25008+c26008+c27008+c28008+c29008+c2A008+c2B008+c2C008+c2D008+c2E008+c2F008;
assign A2008=(C2008>=0)?1:0;

assign P3008=A2008;

ninexnine_unit ninexnine_unit_4132(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20018)
);

ninexnine_unit ninexnine_unit_4133(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21018)
);

ninexnine_unit ninexnine_unit_4134(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22018)
);

ninexnine_unit ninexnine_unit_4135(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23018)
);

ninexnine_unit ninexnine_unit_4136(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24018)
);

ninexnine_unit ninexnine_unit_4137(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25018)
);

ninexnine_unit ninexnine_unit_4138(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26018)
);

ninexnine_unit ninexnine_unit_4139(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27018)
);

ninexnine_unit ninexnine_unit_4140(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W28008),
				.b1(W28018),
				.b2(W28028),
				.b3(W28108),
				.b4(W28118),
				.b5(W28128),
				.b6(W28208),
				.b7(W28218),
				.b8(W28228),
				.c(c28018)
);

ninexnine_unit ninexnine_unit_4141(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W28009),
				.b1(W28019),
				.b2(W28029),
				.b3(W28109),
				.b4(W28119),
				.b5(W28129),
				.b6(W28209),
				.b7(W28219),
				.b8(W28229),
				.c(c29018)
);

ninexnine_unit ninexnine_unit_4142(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2800A),
				.b1(W2801A),
				.b2(W2802A),
				.b3(W2810A),
				.b4(W2811A),
				.b5(W2812A),
				.b6(W2820A),
				.b7(W2821A),
				.b8(W2822A),
				.c(c2A018)
);

ninexnine_unit ninexnine_unit_4143(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2800B),
				.b1(W2801B),
				.b2(W2802B),
				.b3(W2810B),
				.b4(W2811B),
				.b5(W2812B),
				.b6(W2820B),
				.b7(W2821B),
				.b8(W2822B),
				.c(c2B018)
);

ninexnine_unit ninexnine_unit_4144(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2800C),
				.b1(W2801C),
				.b2(W2802C),
				.b3(W2810C),
				.b4(W2811C),
				.b5(W2812C),
				.b6(W2820C),
				.b7(W2821C),
				.b8(W2822C),
				.c(c2C018)
);

ninexnine_unit ninexnine_unit_4145(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2800D),
				.b1(W2801D),
				.b2(W2802D),
				.b3(W2810D),
				.b4(W2811D),
				.b5(W2812D),
				.b6(W2820D),
				.b7(W2821D),
				.b8(W2822D),
				.c(c2D018)
);

ninexnine_unit ninexnine_unit_4146(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2800E),
				.b1(W2801E),
				.b2(W2802E),
				.b3(W2810E),
				.b4(W2811E),
				.b5(W2812E),
				.b6(W2820E),
				.b7(W2821E),
				.b8(W2822E),
				.c(c2E018)
);

ninexnine_unit ninexnine_unit_4147(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2800F),
				.b1(W2801F),
				.b2(W2802F),
				.b3(W2810F),
				.b4(W2811F),
				.b5(W2812F),
				.b6(W2820F),
				.b7(W2821F),
				.b8(W2822F),
				.c(c2F018)
);

assign C2018=c20018+c21018+c22018+c23018+c24018+c25018+c26018+c27018+c28018+c29018+c2A018+c2B018+c2C018+c2D018+c2E018+c2F018;
assign A2018=(C2018>=0)?1:0;

assign P3018=A2018;

ninexnine_unit ninexnine_unit_4148(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20028)
);

ninexnine_unit ninexnine_unit_4149(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21028)
);

ninexnine_unit ninexnine_unit_4150(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22028)
);

ninexnine_unit ninexnine_unit_4151(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23028)
);

ninexnine_unit ninexnine_unit_4152(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24028)
);

ninexnine_unit ninexnine_unit_4153(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25028)
);

ninexnine_unit ninexnine_unit_4154(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26028)
);

ninexnine_unit ninexnine_unit_4155(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27028)
);

ninexnine_unit ninexnine_unit_4156(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W28008),
				.b1(W28018),
				.b2(W28028),
				.b3(W28108),
				.b4(W28118),
				.b5(W28128),
				.b6(W28208),
				.b7(W28218),
				.b8(W28228),
				.c(c28028)
);

ninexnine_unit ninexnine_unit_4157(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W28009),
				.b1(W28019),
				.b2(W28029),
				.b3(W28109),
				.b4(W28119),
				.b5(W28129),
				.b6(W28209),
				.b7(W28219),
				.b8(W28229),
				.c(c29028)
);

ninexnine_unit ninexnine_unit_4158(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2800A),
				.b1(W2801A),
				.b2(W2802A),
				.b3(W2810A),
				.b4(W2811A),
				.b5(W2812A),
				.b6(W2820A),
				.b7(W2821A),
				.b8(W2822A),
				.c(c2A028)
);

ninexnine_unit ninexnine_unit_4159(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2800B),
				.b1(W2801B),
				.b2(W2802B),
				.b3(W2810B),
				.b4(W2811B),
				.b5(W2812B),
				.b6(W2820B),
				.b7(W2821B),
				.b8(W2822B),
				.c(c2B028)
);

ninexnine_unit ninexnine_unit_4160(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2800C),
				.b1(W2801C),
				.b2(W2802C),
				.b3(W2810C),
				.b4(W2811C),
				.b5(W2812C),
				.b6(W2820C),
				.b7(W2821C),
				.b8(W2822C),
				.c(c2C028)
);

ninexnine_unit ninexnine_unit_4161(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2800D),
				.b1(W2801D),
				.b2(W2802D),
				.b3(W2810D),
				.b4(W2811D),
				.b5(W2812D),
				.b6(W2820D),
				.b7(W2821D),
				.b8(W2822D),
				.c(c2D028)
);

ninexnine_unit ninexnine_unit_4162(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2800E),
				.b1(W2801E),
				.b2(W2802E),
				.b3(W2810E),
				.b4(W2811E),
				.b5(W2812E),
				.b6(W2820E),
				.b7(W2821E),
				.b8(W2822E),
				.c(c2E028)
);

ninexnine_unit ninexnine_unit_4163(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2800F),
				.b1(W2801F),
				.b2(W2802F),
				.b3(W2810F),
				.b4(W2811F),
				.b5(W2812F),
				.b6(W2820F),
				.b7(W2821F),
				.b8(W2822F),
				.c(c2F028)
);

assign C2028=c20028+c21028+c22028+c23028+c24028+c25028+c26028+c27028+c28028+c29028+c2A028+c2B028+c2C028+c2D028+c2E028+c2F028;
assign A2028=(C2028>=0)?1:0;

assign P3028=A2028;

ninexnine_unit ninexnine_unit_4164(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20108)
);

ninexnine_unit ninexnine_unit_4165(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21108)
);

ninexnine_unit ninexnine_unit_4166(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22108)
);

ninexnine_unit ninexnine_unit_4167(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23108)
);

ninexnine_unit ninexnine_unit_4168(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24108)
);

ninexnine_unit ninexnine_unit_4169(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25108)
);

ninexnine_unit ninexnine_unit_4170(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26108)
);

ninexnine_unit ninexnine_unit_4171(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27108)
);

ninexnine_unit ninexnine_unit_4172(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W28008),
				.b1(W28018),
				.b2(W28028),
				.b3(W28108),
				.b4(W28118),
				.b5(W28128),
				.b6(W28208),
				.b7(W28218),
				.b8(W28228),
				.c(c28108)
);

ninexnine_unit ninexnine_unit_4173(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W28009),
				.b1(W28019),
				.b2(W28029),
				.b3(W28109),
				.b4(W28119),
				.b5(W28129),
				.b6(W28209),
				.b7(W28219),
				.b8(W28229),
				.c(c29108)
);

ninexnine_unit ninexnine_unit_4174(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2800A),
				.b1(W2801A),
				.b2(W2802A),
				.b3(W2810A),
				.b4(W2811A),
				.b5(W2812A),
				.b6(W2820A),
				.b7(W2821A),
				.b8(W2822A),
				.c(c2A108)
);

ninexnine_unit ninexnine_unit_4175(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2800B),
				.b1(W2801B),
				.b2(W2802B),
				.b3(W2810B),
				.b4(W2811B),
				.b5(W2812B),
				.b6(W2820B),
				.b7(W2821B),
				.b8(W2822B),
				.c(c2B108)
);

ninexnine_unit ninexnine_unit_4176(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2800C),
				.b1(W2801C),
				.b2(W2802C),
				.b3(W2810C),
				.b4(W2811C),
				.b5(W2812C),
				.b6(W2820C),
				.b7(W2821C),
				.b8(W2822C),
				.c(c2C108)
);

ninexnine_unit ninexnine_unit_4177(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2800D),
				.b1(W2801D),
				.b2(W2802D),
				.b3(W2810D),
				.b4(W2811D),
				.b5(W2812D),
				.b6(W2820D),
				.b7(W2821D),
				.b8(W2822D),
				.c(c2D108)
);

ninexnine_unit ninexnine_unit_4178(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2800E),
				.b1(W2801E),
				.b2(W2802E),
				.b3(W2810E),
				.b4(W2811E),
				.b5(W2812E),
				.b6(W2820E),
				.b7(W2821E),
				.b8(W2822E),
				.c(c2E108)
);

ninexnine_unit ninexnine_unit_4179(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2800F),
				.b1(W2801F),
				.b2(W2802F),
				.b3(W2810F),
				.b4(W2811F),
				.b5(W2812F),
				.b6(W2820F),
				.b7(W2821F),
				.b8(W2822F),
				.c(c2F108)
);

assign C2108=c20108+c21108+c22108+c23108+c24108+c25108+c26108+c27108+c28108+c29108+c2A108+c2B108+c2C108+c2D108+c2E108+c2F108;
assign A2108=(C2108>=0)?1:0;

assign P3108=A2108;

ninexnine_unit ninexnine_unit_4180(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20118)
);

ninexnine_unit ninexnine_unit_4181(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21118)
);

ninexnine_unit ninexnine_unit_4182(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22118)
);

ninexnine_unit ninexnine_unit_4183(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23118)
);

ninexnine_unit ninexnine_unit_4184(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24118)
);

ninexnine_unit ninexnine_unit_4185(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25118)
);

ninexnine_unit ninexnine_unit_4186(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26118)
);

ninexnine_unit ninexnine_unit_4187(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27118)
);

ninexnine_unit ninexnine_unit_4188(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W28008),
				.b1(W28018),
				.b2(W28028),
				.b3(W28108),
				.b4(W28118),
				.b5(W28128),
				.b6(W28208),
				.b7(W28218),
				.b8(W28228),
				.c(c28118)
);

ninexnine_unit ninexnine_unit_4189(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W28009),
				.b1(W28019),
				.b2(W28029),
				.b3(W28109),
				.b4(W28119),
				.b5(W28129),
				.b6(W28209),
				.b7(W28219),
				.b8(W28229),
				.c(c29118)
);

ninexnine_unit ninexnine_unit_4190(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2800A),
				.b1(W2801A),
				.b2(W2802A),
				.b3(W2810A),
				.b4(W2811A),
				.b5(W2812A),
				.b6(W2820A),
				.b7(W2821A),
				.b8(W2822A),
				.c(c2A118)
);

ninexnine_unit ninexnine_unit_4191(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2800B),
				.b1(W2801B),
				.b2(W2802B),
				.b3(W2810B),
				.b4(W2811B),
				.b5(W2812B),
				.b6(W2820B),
				.b7(W2821B),
				.b8(W2822B),
				.c(c2B118)
);

ninexnine_unit ninexnine_unit_4192(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2800C),
				.b1(W2801C),
				.b2(W2802C),
				.b3(W2810C),
				.b4(W2811C),
				.b5(W2812C),
				.b6(W2820C),
				.b7(W2821C),
				.b8(W2822C),
				.c(c2C118)
);

ninexnine_unit ninexnine_unit_4193(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2800D),
				.b1(W2801D),
				.b2(W2802D),
				.b3(W2810D),
				.b4(W2811D),
				.b5(W2812D),
				.b6(W2820D),
				.b7(W2821D),
				.b8(W2822D),
				.c(c2D118)
);

ninexnine_unit ninexnine_unit_4194(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2800E),
				.b1(W2801E),
				.b2(W2802E),
				.b3(W2810E),
				.b4(W2811E),
				.b5(W2812E),
				.b6(W2820E),
				.b7(W2821E),
				.b8(W2822E),
				.c(c2E118)
);

ninexnine_unit ninexnine_unit_4195(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2800F),
				.b1(W2801F),
				.b2(W2802F),
				.b3(W2810F),
				.b4(W2811F),
				.b5(W2812F),
				.b6(W2820F),
				.b7(W2821F),
				.b8(W2822F),
				.c(c2F118)
);

assign C2118=c20118+c21118+c22118+c23118+c24118+c25118+c26118+c27118+c28118+c29118+c2A118+c2B118+c2C118+c2D118+c2E118+c2F118;
assign A2118=(C2118>=0)?1:0;

assign P3118=A2118;

ninexnine_unit ninexnine_unit_4196(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20128)
);

ninexnine_unit ninexnine_unit_4197(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21128)
);

ninexnine_unit ninexnine_unit_4198(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22128)
);

ninexnine_unit ninexnine_unit_4199(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23128)
);

ninexnine_unit ninexnine_unit_4200(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24128)
);

ninexnine_unit ninexnine_unit_4201(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25128)
);

ninexnine_unit ninexnine_unit_4202(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26128)
);

ninexnine_unit ninexnine_unit_4203(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27128)
);

ninexnine_unit ninexnine_unit_4204(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W28008),
				.b1(W28018),
				.b2(W28028),
				.b3(W28108),
				.b4(W28118),
				.b5(W28128),
				.b6(W28208),
				.b7(W28218),
				.b8(W28228),
				.c(c28128)
);

ninexnine_unit ninexnine_unit_4205(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W28009),
				.b1(W28019),
				.b2(W28029),
				.b3(W28109),
				.b4(W28119),
				.b5(W28129),
				.b6(W28209),
				.b7(W28219),
				.b8(W28229),
				.c(c29128)
);

ninexnine_unit ninexnine_unit_4206(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2800A),
				.b1(W2801A),
				.b2(W2802A),
				.b3(W2810A),
				.b4(W2811A),
				.b5(W2812A),
				.b6(W2820A),
				.b7(W2821A),
				.b8(W2822A),
				.c(c2A128)
);

ninexnine_unit ninexnine_unit_4207(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2800B),
				.b1(W2801B),
				.b2(W2802B),
				.b3(W2810B),
				.b4(W2811B),
				.b5(W2812B),
				.b6(W2820B),
				.b7(W2821B),
				.b8(W2822B),
				.c(c2B128)
);

ninexnine_unit ninexnine_unit_4208(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2800C),
				.b1(W2801C),
				.b2(W2802C),
				.b3(W2810C),
				.b4(W2811C),
				.b5(W2812C),
				.b6(W2820C),
				.b7(W2821C),
				.b8(W2822C),
				.c(c2C128)
);

ninexnine_unit ninexnine_unit_4209(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2800D),
				.b1(W2801D),
				.b2(W2802D),
				.b3(W2810D),
				.b4(W2811D),
				.b5(W2812D),
				.b6(W2820D),
				.b7(W2821D),
				.b8(W2822D),
				.c(c2D128)
);

ninexnine_unit ninexnine_unit_4210(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2800E),
				.b1(W2801E),
				.b2(W2802E),
				.b3(W2810E),
				.b4(W2811E),
				.b5(W2812E),
				.b6(W2820E),
				.b7(W2821E),
				.b8(W2822E),
				.c(c2E128)
);

ninexnine_unit ninexnine_unit_4211(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2800F),
				.b1(W2801F),
				.b2(W2802F),
				.b3(W2810F),
				.b4(W2811F),
				.b5(W2812F),
				.b6(W2820F),
				.b7(W2821F),
				.b8(W2822F),
				.c(c2F128)
);

assign C2128=c20128+c21128+c22128+c23128+c24128+c25128+c26128+c27128+c28128+c29128+c2A128+c2B128+c2C128+c2D128+c2E128+c2F128;
assign A2128=(C2128>=0)?1:0;

assign P3128=A2128;

ninexnine_unit ninexnine_unit_4212(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20208)
);

ninexnine_unit ninexnine_unit_4213(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21208)
);

ninexnine_unit ninexnine_unit_4214(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22208)
);

ninexnine_unit ninexnine_unit_4215(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23208)
);

ninexnine_unit ninexnine_unit_4216(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24208)
);

ninexnine_unit ninexnine_unit_4217(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25208)
);

ninexnine_unit ninexnine_unit_4218(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26208)
);

ninexnine_unit ninexnine_unit_4219(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27208)
);

ninexnine_unit ninexnine_unit_4220(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W28008),
				.b1(W28018),
				.b2(W28028),
				.b3(W28108),
				.b4(W28118),
				.b5(W28128),
				.b6(W28208),
				.b7(W28218),
				.b8(W28228),
				.c(c28208)
);

ninexnine_unit ninexnine_unit_4221(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W28009),
				.b1(W28019),
				.b2(W28029),
				.b3(W28109),
				.b4(W28119),
				.b5(W28129),
				.b6(W28209),
				.b7(W28219),
				.b8(W28229),
				.c(c29208)
);

ninexnine_unit ninexnine_unit_4222(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2800A),
				.b1(W2801A),
				.b2(W2802A),
				.b3(W2810A),
				.b4(W2811A),
				.b5(W2812A),
				.b6(W2820A),
				.b7(W2821A),
				.b8(W2822A),
				.c(c2A208)
);

ninexnine_unit ninexnine_unit_4223(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2800B),
				.b1(W2801B),
				.b2(W2802B),
				.b3(W2810B),
				.b4(W2811B),
				.b5(W2812B),
				.b6(W2820B),
				.b7(W2821B),
				.b8(W2822B),
				.c(c2B208)
);

ninexnine_unit ninexnine_unit_4224(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2800C),
				.b1(W2801C),
				.b2(W2802C),
				.b3(W2810C),
				.b4(W2811C),
				.b5(W2812C),
				.b6(W2820C),
				.b7(W2821C),
				.b8(W2822C),
				.c(c2C208)
);

ninexnine_unit ninexnine_unit_4225(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2800D),
				.b1(W2801D),
				.b2(W2802D),
				.b3(W2810D),
				.b4(W2811D),
				.b5(W2812D),
				.b6(W2820D),
				.b7(W2821D),
				.b8(W2822D),
				.c(c2D208)
);

ninexnine_unit ninexnine_unit_4226(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2800E),
				.b1(W2801E),
				.b2(W2802E),
				.b3(W2810E),
				.b4(W2811E),
				.b5(W2812E),
				.b6(W2820E),
				.b7(W2821E),
				.b8(W2822E),
				.c(c2E208)
);

ninexnine_unit ninexnine_unit_4227(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2800F),
				.b1(W2801F),
				.b2(W2802F),
				.b3(W2810F),
				.b4(W2811F),
				.b5(W2812F),
				.b6(W2820F),
				.b7(W2821F),
				.b8(W2822F),
				.c(c2F208)
);

assign C2208=c20208+c21208+c22208+c23208+c24208+c25208+c26208+c27208+c28208+c29208+c2A208+c2B208+c2C208+c2D208+c2E208+c2F208;
assign A2208=(C2208>=0)?1:0;

assign P3208=A2208;

ninexnine_unit ninexnine_unit_4228(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20218)
);

ninexnine_unit ninexnine_unit_4229(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21218)
);

ninexnine_unit ninexnine_unit_4230(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22218)
);

ninexnine_unit ninexnine_unit_4231(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23218)
);

ninexnine_unit ninexnine_unit_4232(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24218)
);

ninexnine_unit ninexnine_unit_4233(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25218)
);

ninexnine_unit ninexnine_unit_4234(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26218)
);

ninexnine_unit ninexnine_unit_4235(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27218)
);

ninexnine_unit ninexnine_unit_4236(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W28008),
				.b1(W28018),
				.b2(W28028),
				.b3(W28108),
				.b4(W28118),
				.b5(W28128),
				.b6(W28208),
				.b7(W28218),
				.b8(W28228),
				.c(c28218)
);

ninexnine_unit ninexnine_unit_4237(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W28009),
				.b1(W28019),
				.b2(W28029),
				.b3(W28109),
				.b4(W28119),
				.b5(W28129),
				.b6(W28209),
				.b7(W28219),
				.b8(W28229),
				.c(c29218)
);

ninexnine_unit ninexnine_unit_4238(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2800A),
				.b1(W2801A),
				.b2(W2802A),
				.b3(W2810A),
				.b4(W2811A),
				.b5(W2812A),
				.b6(W2820A),
				.b7(W2821A),
				.b8(W2822A),
				.c(c2A218)
);

ninexnine_unit ninexnine_unit_4239(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2800B),
				.b1(W2801B),
				.b2(W2802B),
				.b3(W2810B),
				.b4(W2811B),
				.b5(W2812B),
				.b6(W2820B),
				.b7(W2821B),
				.b8(W2822B),
				.c(c2B218)
);

ninexnine_unit ninexnine_unit_4240(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2800C),
				.b1(W2801C),
				.b2(W2802C),
				.b3(W2810C),
				.b4(W2811C),
				.b5(W2812C),
				.b6(W2820C),
				.b7(W2821C),
				.b8(W2822C),
				.c(c2C218)
);

ninexnine_unit ninexnine_unit_4241(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2800D),
				.b1(W2801D),
				.b2(W2802D),
				.b3(W2810D),
				.b4(W2811D),
				.b5(W2812D),
				.b6(W2820D),
				.b7(W2821D),
				.b8(W2822D),
				.c(c2D218)
);

ninexnine_unit ninexnine_unit_4242(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2800E),
				.b1(W2801E),
				.b2(W2802E),
				.b3(W2810E),
				.b4(W2811E),
				.b5(W2812E),
				.b6(W2820E),
				.b7(W2821E),
				.b8(W2822E),
				.c(c2E218)
);

ninexnine_unit ninexnine_unit_4243(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2800F),
				.b1(W2801F),
				.b2(W2802F),
				.b3(W2810F),
				.b4(W2811F),
				.b5(W2812F),
				.b6(W2820F),
				.b7(W2821F),
				.b8(W2822F),
				.c(c2F218)
);

assign C2218=c20218+c21218+c22218+c23218+c24218+c25218+c26218+c27218+c28218+c29218+c2A218+c2B218+c2C218+c2D218+c2E218+c2F218;
assign A2218=(C2218>=0)?1:0;

assign P3218=A2218;

ninexnine_unit ninexnine_unit_4244(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W28000),
				.b1(W28010),
				.b2(W28020),
				.b3(W28100),
				.b4(W28110),
				.b5(W28120),
				.b6(W28200),
				.b7(W28210),
				.b8(W28220),
				.c(c20228)
);

ninexnine_unit ninexnine_unit_4245(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W28001),
				.b1(W28011),
				.b2(W28021),
				.b3(W28101),
				.b4(W28111),
				.b5(W28121),
				.b6(W28201),
				.b7(W28211),
				.b8(W28221),
				.c(c21228)
);

ninexnine_unit ninexnine_unit_4246(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W28002),
				.b1(W28012),
				.b2(W28022),
				.b3(W28102),
				.b4(W28112),
				.b5(W28122),
				.b6(W28202),
				.b7(W28212),
				.b8(W28222),
				.c(c22228)
);

ninexnine_unit ninexnine_unit_4247(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W28003),
				.b1(W28013),
				.b2(W28023),
				.b3(W28103),
				.b4(W28113),
				.b5(W28123),
				.b6(W28203),
				.b7(W28213),
				.b8(W28223),
				.c(c23228)
);

ninexnine_unit ninexnine_unit_4248(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W28004),
				.b1(W28014),
				.b2(W28024),
				.b3(W28104),
				.b4(W28114),
				.b5(W28124),
				.b6(W28204),
				.b7(W28214),
				.b8(W28224),
				.c(c24228)
);

ninexnine_unit ninexnine_unit_4249(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W28005),
				.b1(W28015),
				.b2(W28025),
				.b3(W28105),
				.b4(W28115),
				.b5(W28125),
				.b6(W28205),
				.b7(W28215),
				.b8(W28225),
				.c(c25228)
);

ninexnine_unit ninexnine_unit_4250(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W28006),
				.b1(W28016),
				.b2(W28026),
				.b3(W28106),
				.b4(W28116),
				.b5(W28126),
				.b6(W28206),
				.b7(W28216),
				.b8(W28226),
				.c(c26228)
);

ninexnine_unit ninexnine_unit_4251(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W28007),
				.b1(W28017),
				.b2(W28027),
				.b3(W28107),
				.b4(W28117),
				.b5(W28127),
				.b6(W28207),
				.b7(W28217),
				.b8(W28227),
				.c(c27228)
);

ninexnine_unit ninexnine_unit_4252(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W28008),
				.b1(W28018),
				.b2(W28028),
				.b3(W28108),
				.b4(W28118),
				.b5(W28128),
				.b6(W28208),
				.b7(W28218),
				.b8(W28228),
				.c(c28228)
);

ninexnine_unit ninexnine_unit_4253(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W28009),
				.b1(W28019),
				.b2(W28029),
				.b3(W28109),
				.b4(W28119),
				.b5(W28129),
				.b6(W28209),
				.b7(W28219),
				.b8(W28229),
				.c(c29228)
);

ninexnine_unit ninexnine_unit_4254(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2800A),
				.b1(W2801A),
				.b2(W2802A),
				.b3(W2810A),
				.b4(W2811A),
				.b5(W2812A),
				.b6(W2820A),
				.b7(W2821A),
				.b8(W2822A),
				.c(c2A228)
);

ninexnine_unit ninexnine_unit_4255(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2800B),
				.b1(W2801B),
				.b2(W2802B),
				.b3(W2810B),
				.b4(W2811B),
				.b5(W2812B),
				.b6(W2820B),
				.b7(W2821B),
				.b8(W2822B),
				.c(c2B228)
);

ninexnine_unit ninexnine_unit_4256(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2800C),
				.b1(W2801C),
				.b2(W2802C),
				.b3(W2810C),
				.b4(W2811C),
				.b5(W2812C),
				.b6(W2820C),
				.b7(W2821C),
				.b8(W2822C),
				.c(c2C228)
);

ninexnine_unit ninexnine_unit_4257(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2800D),
				.b1(W2801D),
				.b2(W2802D),
				.b3(W2810D),
				.b4(W2811D),
				.b5(W2812D),
				.b6(W2820D),
				.b7(W2821D),
				.b8(W2822D),
				.c(c2D228)
);

ninexnine_unit ninexnine_unit_4258(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2800E),
				.b1(W2801E),
				.b2(W2802E),
				.b3(W2810E),
				.b4(W2811E),
				.b5(W2812E),
				.b6(W2820E),
				.b7(W2821E),
				.b8(W2822E),
				.c(c2E228)
);

ninexnine_unit ninexnine_unit_4259(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2800F),
				.b1(W2801F),
				.b2(W2802F),
				.b3(W2810F),
				.b4(W2811F),
				.b5(W2812F),
				.b6(W2820F),
				.b7(W2821F),
				.b8(W2822F),
				.c(c2F228)
);

assign C2228=c20228+c21228+c22228+c23228+c24228+c25228+c26228+c27228+c28228+c29228+c2A228+c2B228+c2C228+c2D228+c2E228+c2F228;
assign A2228=(C2228>=0)?1:0;

assign P3228=A2228;

ninexnine_unit ninexnine_unit_4260(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20009)
);

ninexnine_unit ninexnine_unit_4261(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21009)
);

ninexnine_unit ninexnine_unit_4262(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22009)
);

ninexnine_unit ninexnine_unit_4263(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23009)
);

ninexnine_unit ninexnine_unit_4264(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24009)
);

ninexnine_unit ninexnine_unit_4265(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25009)
);

ninexnine_unit ninexnine_unit_4266(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26009)
);

ninexnine_unit ninexnine_unit_4267(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27009)
);

ninexnine_unit ninexnine_unit_4268(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W29008),
				.b1(W29018),
				.b2(W29028),
				.b3(W29108),
				.b4(W29118),
				.b5(W29128),
				.b6(W29208),
				.b7(W29218),
				.b8(W29228),
				.c(c28009)
);

ninexnine_unit ninexnine_unit_4269(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W29009),
				.b1(W29019),
				.b2(W29029),
				.b3(W29109),
				.b4(W29119),
				.b5(W29129),
				.b6(W29209),
				.b7(W29219),
				.b8(W29229),
				.c(c29009)
);

ninexnine_unit ninexnine_unit_4270(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2900A),
				.b1(W2901A),
				.b2(W2902A),
				.b3(W2910A),
				.b4(W2911A),
				.b5(W2912A),
				.b6(W2920A),
				.b7(W2921A),
				.b8(W2922A),
				.c(c2A009)
);

ninexnine_unit ninexnine_unit_4271(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2900B),
				.b1(W2901B),
				.b2(W2902B),
				.b3(W2910B),
				.b4(W2911B),
				.b5(W2912B),
				.b6(W2920B),
				.b7(W2921B),
				.b8(W2922B),
				.c(c2B009)
);

ninexnine_unit ninexnine_unit_4272(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2900C),
				.b1(W2901C),
				.b2(W2902C),
				.b3(W2910C),
				.b4(W2911C),
				.b5(W2912C),
				.b6(W2920C),
				.b7(W2921C),
				.b8(W2922C),
				.c(c2C009)
);

ninexnine_unit ninexnine_unit_4273(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2900D),
				.b1(W2901D),
				.b2(W2902D),
				.b3(W2910D),
				.b4(W2911D),
				.b5(W2912D),
				.b6(W2920D),
				.b7(W2921D),
				.b8(W2922D),
				.c(c2D009)
);

ninexnine_unit ninexnine_unit_4274(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2900E),
				.b1(W2901E),
				.b2(W2902E),
				.b3(W2910E),
				.b4(W2911E),
				.b5(W2912E),
				.b6(W2920E),
				.b7(W2921E),
				.b8(W2922E),
				.c(c2E009)
);

ninexnine_unit ninexnine_unit_4275(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2900F),
				.b1(W2901F),
				.b2(W2902F),
				.b3(W2910F),
				.b4(W2911F),
				.b5(W2912F),
				.b6(W2920F),
				.b7(W2921F),
				.b8(W2922F),
				.c(c2F009)
);

assign C2009=c20009+c21009+c22009+c23009+c24009+c25009+c26009+c27009+c28009+c29009+c2A009+c2B009+c2C009+c2D009+c2E009+c2F009;
assign A2009=(C2009>=0)?1:0;

assign P3009=A2009;

ninexnine_unit ninexnine_unit_4276(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20019)
);

ninexnine_unit ninexnine_unit_4277(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21019)
);

ninexnine_unit ninexnine_unit_4278(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22019)
);

ninexnine_unit ninexnine_unit_4279(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23019)
);

ninexnine_unit ninexnine_unit_4280(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24019)
);

ninexnine_unit ninexnine_unit_4281(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25019)
);

ninexnine_unit ninexnine_unit_4282(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26019)
);

ninexnine_unit ninexnine_unit_4283(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27019)
);

ninexnine_unit ninexnine_unit_4284(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W29008),
				.b1(W29018),
				.b2(W29028),
				.b3(W29108),
				.b4(W29118),
				.b5(W29128),
				.b6(W29208),
				.b7(W29218),
				.b8(W29228),
				.c(c28019)
);

ninexnine_unit ninexnine_unit_4285(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W29009),
				.b1(W29019),
				.b2(W29029),
				.b3(W29109),
				.b4(W29119),
				.b5(W29129),
				.b6(W29209),
				.b7(W29219),
				.b8(W29229),
				.c(c29019)
);

ninexnine_unit ninexnine_unit_4286(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2900A),
				.b1(W2901A),
				.b2(W2902A),
				.b3(W2910A),
				.b4(W2911A),
				.b5(W2912A),
				.b6(W2920A),
				.b7(W2921A),
				.b8(W2922A),
				.c(c2A019)
);

ninexnine_unit ninexnine_unit_4287(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2900B),
				.b1(W2901B),
				.b2(W2902B),
				.b3(W2910B),
				.b4(W2911B),
				.b5(W2912B),
				.b6(W2920B),
				.b7(W2921B),
				.b8(W2922B),
				.c(c2B019)
);

ninexnine_unit ninexnine_unit_4288(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2900C),
				.b1(W2901C),
				.b2(W2902C),
				.b3(W2910C),
				.b4(W2911C),
				.b5(W2912C),
				.b6(W2920C),
				.b7(W2921C),
				.b8(W2922C),
				.c(c2C019)
);

ninexnine_unit ninexnine_unit_4289(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2900D),
				.b1(W2901D),
				.b2(W2902D),
				.b3(W2910D),
				.b4(W2911D),
				.b5(W2912D),
				.b6(W2920D),
				.b7(W2921D),
				.b8(W2922D),
				.c(c2D019)
);

ninexnine_unit ninexnine_unit_4290(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2900E),
				.b1(W2901E),
				.b2(W2902E),
				.b3(W2910E),
				.b4(W2911E),
				.b5(W2912E),
				.b6(W2920E),
				.b7(W2921E),
				.b8(W2922E),
				.c(c2E019)
);

ninexnine_unit ninexnine_unit_4291(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2900F),
				.b1(W2901F),
				.b2(W2902F),
				.b3(W2910F),
				.b4(W2911F),
				.b5(W2912F),
				.b6(W2920F),
				.b7(W2921F),
				.b8(W2922F),
				.c(c2F019)
);

assign C2019=c20019+c21019+c22019+c23019+c24019+c25019+c26019+c27019+c28019+c29019+c2A019+c2B019+c2C019+c2D019+c2E019+c2F019;
assign A2019=(C2019>=0)?1:0;

assign P3019=A2019;

ninexnine_unit ninexnine_unit_4292(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20029)
);

ninexnine_unit ninexnine_unit_4293(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21029)
);

ninexnine_unit ninexnine_unit_4294(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22029)
);

ninexnine_unit ninexnine_unit_4295(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23029)
);

ninexnine_unit ninexnine_unit_4296(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24029)
);

ninexnine_unit ninexnine_unit_4297(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25029)
);

ninexnine_unit ninexnine_unit_4298(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26029)
);

ninexnine_unit ninexnine_unit_4299(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27029)
);

ninexnine_unit ninexnine_unit_4300(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W29008),
				.b1(W29018),
				.b2(W29028),
				.b3(W29108),
				.b4(W29118),
				.b5(W29128),
				.b6(W29208),
				.b7(W29218),
				.b8(W29228),
				.c(c28029)
);

ninexnine_unit ninexnine_unit_4301(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W29009),
				.b1(W29019),
				.b2(W29029),
				.b3(W29109),
				.b4(W29119),
				.b5(W29129),
				.b6(W29209),
				.b7(W29219),
				.b8(W29229),
				.c(c29029)
);

ninexnine_unit ninexnine_unit_4302(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2900A),
				.b1(W2901A),
				.b2(W2902A),
				.b3(W2910A),
				.b4(W2911A),
				.b5(W2912A),
				.b6(W2920A),
				.b7(W2921A),
				.b8(W2922A),
				.c(c2A029)
);

ninexnine_unit ninexnine_unit_4303(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2900B),
				.b1(W2901B),
				.b2(W2902B),
				.b3(W2910B),
				.b4(W2911B),
				.b5(W2912B),
				.b6(W2920B),
				.b7(W2921B),
				.b8(W2922B),
				.c(c2B029)
);

ninexnine_unit ninexnine_unit_4304(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2900C),
				.b1(W2901C),
				.b2(W2902C),
				.b3(W2910C),
				.b4(W2911C),
				.b5(W2912C),
				.b6(W2920C),
				.b7(W2921C),
				.b8(W2922C),
				.c(c2C029)
);

ninexnine_unit ninexnine_unit_4305(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2900D),
				.b1(W2901D),
				.b2(W2902D),
				.b3(W2910D),
				.b4(W2911D),
				.b5(W2912D),
				.b6(W2920D),
				.b7(W2921D),
				.b8(W2922D),
				.c(c2D029)
);

ninexnine_unit ninexnine_unit_4306(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2900E),
				.b1(W2901E),
				.b2(W2902E),
				.b3(W2910E),
				.b4(W2911E),
				.b5(W2912E),
				.b6(W2920E),
				.b7(W2921E),
				.b8(W2922E),
				.c(c2E029)
);

ninexnine_unit ninexnine_unit_4307(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2900F),
				.b1(W2901F),
				.b2(W2902F),
				.b3(W2910F),
				.b4(W2911F),
				.b5(W2912F),
				.b6(W2920F),
				.b7(W2921F),
				.b8(W2922F),
				.c(c2F029)
);

assign C2029=c20029+c21029+c22029+c23029+c24029+c25029+c26029+c27029+c28029+c29029+c2A029+c2B029+c2C029+c2D029+c2E029+c2F029;
assign A2029=(C2029>=0)?1:0;

assign P3029=A2029;

ninexnine_unit ninexnine_unit_4308(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20109)
);

ninexnine_unit ninexnine_unit_4309(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21109)
);

ninexnine_unit ninexnine_unit_4310(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22109)
);

ninexnine_unit ninexnine_unit_4311(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23109)
);

ninexnine_unit ninexnine_unit_4312(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24109)
);

ninexnine_unit ninexnine_unit_4313(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25109)
);

ninexnine_unit ninexnine_unit_4314(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26109)
);

ninexnine_unit ninexnine_unit_4315(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27109)
);

ninexnine_unit ninexnine_unit_4316(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W29008),
				.b1(W29018),
				.b2(W29028),
				.b3(W29108),
				.b4(W29118),
				.b5(W29128),
				.b6(W29208),
				.b7(W29218),
				.b8(W29228),
				.c(c28109)
);

ninexnine_unit ninexnine_unit_4317(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W29009),
				.b1(W29019),
				.b2(W29029),
				.b3(W29109),
				.b4(W29119),
				.b5(W29129),
				.b6(W29209),
				.b7(W29219),
				.b8(W29229),
				.c(c29109)
);

ninexnine_unit ninexnine_unit_4318(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2900A),
				.b1(W2901A),
				.b2(W2902A),
				.b3(W2910A),
				.b4(W2911A),
				.b5(W2912A),
				.b6(W2920A),
				.b7(W2921A),
				.b8(W2922A),
				.c(c2A109)
);

ninexnine_unit ninexnine_unit_4319(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2900B),
				.b1(W2901B),
				.b2(W2902B),
				.b3(W2910B),
				.b4(W2911B),
				.b5(W2912B),
				.b6(W2920B),
				.b7(W2921B),
				.b8(W2922B),
				.c(c2B109)
);

ninexnine_unit ninexnine_unit_4320(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2900C),
				.b1(W2901C),
				.b2(W2902C),
				.b3(W2910C),
				.b4(W2911C),
				.b5(W2912C),
				.b6(W2920C),
				.b7(W2921C),
				.b8(W2922C),
				.c(c2C109)
);

ninexnine_unit ninexnine_unit_4321(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2900D),
				.b1(W2901D),
				.b2(W2902D),
				.b3(W2910D),
				.b4(W2911D),
				.b5(W2912D),
				.b6(W2920D),
				.b7(W2921D),
				.b8(W2922D),
				.c(c2D109)
);

ninexnine_unit ninexnine_unit_4322(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2900E),
				.b1(W2901E),
				.b2(W2902E),
				.b3(W2910E),
				.b4(W2911E),
				.b5(W2912E),
				.b6(W2920E),
				.b7(W2921E),
				.b8(W2922E),
				.c(c2E109)
);

ninexnine_unit ninexnine_unit_4323(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2900F),
				.b1(W2901F),
				.b2(W2902F),
				.b3(W2910F),
				.b4(W2911F),
				.b5(W2912F),
				.b6(W2920F),
				.b7(W2921F),
				.b8(W2922F),
				.c(c2F109)
);

assign C2109=c20109+c21109+c22109+c23109+c24109+c25109+c26109+c27109+c28109+c29109+c2A109+c2B109+c2C109+c2D109+c2E109+c2F109;
assign A2109=(C2109>=0)?1:0;

assign P3109=A2109;

ninexnine_unit ninexnine_unit_4324(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20119)
);

ninexnine_unit ninexnine_unit_4325(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21119)
);

ninexnine_unit ninexnine_unit_4326(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22119)
);

ninexnine_unit ninexnine_unit_4327(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23119)
);

ninexnine_unit ninexnine_unit_4328(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24119)
);

ninexnine_unit ninexnine_unit_4329(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25119)
);

ninexnine_unit ninexnine_unit_4330(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26119)
);

ninexnine_unit ninexnine_unit_4331(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27119)
);

ninexnine_unit ninexnine_unit_4332(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W29008),
				.b1(W29018),
				.b2(W29028),
				.b3(W29108),
				.b4(W29118),
				.b5(W29128),
				.b6(W29208),
				.b7(W29218),
				.b8(W29228),
				.c(c28119)
);

ninexnine_unit ninexnine_unit_4333(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W29009),
				.b1(W29019),
				.b2(W29029),
				.b3(W29109),
				.b4(W29119),
				.b5(W29129),
				.b6(W29209),
				.b7(W29219),
				.b8(W29229),
				.c(c29119)
);

ninexnine_unit ninexnine_unit_4334(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2900A),
				.b1(W2901A),
				.b2(W2902A),
				.b3(W2910A),
				.b4(W2911A),
				.b5(W2912A),
				.b6(W2920A),
				.b7(W2921A),
				.b8(W2922A),
				.c(c2A119)
);

ninexnine_unit ninexnine_unit_4335(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2900B),
				.b1(W2901B),
				.b2(W2902B),
				.b3(W2910B),
				.b4(W2911B),
				.b5(W2912B),
				.b6(W2920B),
				.b7(W2921B),
				.b8(W2922B),
				.c(c2B119)
);

ninexnine_unit ninexnine_unit_4336(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2900C),
				.b1(W2901C),
				.b2(W2902C),
				.b3(W2910C),
				.b4(W2911C),
				.b5(W2912C),
				.b6(W2920C),
				.b7(W2921C),
				.b8(W2922C),
				.c(c2C119)
);

ninexnine_unit ninexnine_unit_4337(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2900D),
				.b1(W2901D),
				.b2(W2902D),
				.b3(W2910D),
				.b4(W2911D),
				.b5(W2912D),
				.b6(W2920D),
				.b7(W2921D),
				.b8(W2922D),
				.c(c2D119)
);

ninexnine_unit ninexnine_unit_4338(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2900E),
				.b1(W2901E),
				.b2(W2902E),
				.b3(W2910E),
				.b4(W2911E),
				.b5(W2912E),
				.b6(W2920E),
				.b7(W2921E),
				.b8(W2922E),
				.c(c2E119)
);

ninexnine_unit ninexnine_unit_4339(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2900F),
				.b1(W2901F),
				.b2(W2902F),
				.b3(W2910F),
				.b4(W2911F),
				.b5(W2912F),
				.b6(W2920F),
				.b7(W2921F),
				.b8(W2922F),
				.c(c2F119)
);

assign C2119=c20119+c21119+c22119+c23119+c24119+c25119+c26119+c27119+c28119+c29119+c2A119+c2B119+c2C119+c2D119+c2E119+c2F119;
assign A2119=(C2119>=0)?1:0;

assign P3119=A2119;

ninexnine_unit ninexnine_unit_4340(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20129)
);

ninexnine_unit ninexnine_unit_4341(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21129)
);

ninexnine_unit ninexnine_unit_4342(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22129)
);

ninexnine_unit ninexnine_unit_4343(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23129)
);

ninexnine_unit ninexnine_unit_4344(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24129)
);

ninexnine_unit ninexnine_unit_4345(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25129)
);

ninexnine_unit ninexnine_unit_4346(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26129)
);

ninexnine_unit ninexnine_unit_4347(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27129)
);

ninexnine_unit ninexnine_unit_4348(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W29008),
				.b1(W29018),
				.b2(W29028),
				.b3(W29108),
				.b4(W29118),
				.b5(W29128),
				.b6(W29208),
				.b7(W29218),
				.b8(W29228),
				.c(c28129)
);

ninexnine_unit ninexnine_unit_4349(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W29009),
				.b1(W29019),
				.b2(W29029),
				.b3(W29109),
				.b4(W29119),
				.b5(W29129),
				.b6(W29209),
				.b7(W29219),
				.b8(W29229),
				.c(c29129)
);

ninexnine_unit ninexnine_unit_4350(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2900A),
				.b1(W2901A),
				.b2(W2902A),
				.b3(W2910A),
				.b4(W2911A),
				.b5(W2912A),
				.b6(W2920A),
				.b7(W2921A),
				.b8(W2922A),
				.c(c2A129)
);

ninexnine_unit ninexnine_unit_4351(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2900B),
				.b1(W2901B),
				.b2(W2902B),
				.b3(W2910B),
				.b4(W2911B),
				.b5(W2912B),
				.b6(W2920B),
				.b7(W2921B),
				.b8(W2922B),
				.c(c2B129)
);

ninexnine_unit ninexnine_unit_4352(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2900C),
				.b1(W2901C),
				.b2(W2902C),
				.b3(W2910C),
				.b4(W2911C),
				.b5(W2912C),
				.b6(W2920C),
				.b7(W2921C),
				.b8(W2922C),
				.c(c2C129)
);

ninexnine_unit ninexnine_unit_4353(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2900D),
				.b1(W2901D),
				.b2(W2902D),
				.b3(W2910D),
				.b4(W2911D),
				.b5(W2912D),
				.b6(W2920D),
				.b7(W2921D),
				.b8(W2922D),
				.c(c2D129)
);

ninexnine_unit ninexnine_unit_4354(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2900E),
				.b1(W2901E),
				.b2(W2902E),
				.b3(W2910E),
				.b4(W2911E),
				.b5(W2912E),
				.b6(W2920E),
				.b7(W2921E),
				.b8(W2922E),
				.c(c2E129)
);

ninexnine_unit ninexnine_unit_4355(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2900F),
				.b1(W2901F),
				.b2(W2902F),
				.b3(W2910F),
				.b4(W2911F),
				.b5(W2912F),
				.b6(W2920F),
				.b7(W2921F),
				.b8(W2922F),
				.c(c2F129)
);

assign C2129=c20129+c21129+c22129+c23129+c24129+c25129+c26129+c27129+c28129+c29129+c2A129+c2B129+c2C129+c2D129+c2E129+c2F129;
assign A2129=(C2129>=0)?1:0;

assign P3129=A2129;

ninexnine_unit ninexnine_unit_4356(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20209)
);

ninexnine_unit ninexnine_unit_4357(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21209)
);

ninexnine_unit ninexnine_unit_4358(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22209)
);

ninexnine_unit ninexnine_unit_4359(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23209)
);

ninexnine_unit ninexnine_unit_4360(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24209)
);

ninexnine_unit ninexnine_unit_4361(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25209)
);

ninexnine_unit ninexnine_unit_4362(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26209)
);

ninexnine_unit ninexnine_unit_4363(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27209)
);

ninexnine_unit ninexnine_unit_4364(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W29008),
				.b1(W29018),
				.b2(W29028),
				.b3(W29108),
				.b4(W29118),
				.b5(W29128),
				.b6(W29208),
				.b7(W29218),
				.b8(W29228),
				.c(c28209)
);

ninexnine_unit ninexnine_unit_4365(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W29009),
				.b1(W29019),
				.b2(W29029),
				.b3(W29109),
				.b4(W29119),
				.b5(W29129),
				.b6(W29209),
				.b7(W29219),
				.b8(W29229),
				.c(c29209)
);

ninexnine_unit ninexnine_unit_4366(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2900A),
				.b1(W2901A),
				.b2(W2902A),
				.b3(W2910A),
				.b4(W2911A),
				.b5(W2912A),
				.b6(W2920A),
				.b7(W2921A),
				.b8(W2922A),
				.c(c2A209)
);

ninexnine_unit ninexnine_unit_4367(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2900B),
				.b1(W2901B),
				.b2(W2902B),
				.b3(W2910B),
				.b4(W2911B),
				.b5(W2912B),
				.b6(W2920B),
				.b7(W2921B),
				.b8(W2922B),
				.c(c2B209)
);

ninexnine_unit ninexnine_unit_4368(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2900C),
				.b1(W2901C),
				.b2(W2902C),
				.b3(W2910C),
				.b4(W2911C),
				.b5(W2912C),
				.b6(W2920C),
				.b7(W2921C),
				.b8(W2922C),
				.c(c2C209)
);

ninexnine_unit ninexnine_unit_4369(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2900D),
				.b1(W2901D),
				.b2(W2902D),
				.b3(W2910D),
				.b4(W2911D),
				.b5(W2912D),
				.b6(W2920D),
				.b7(W2921D),
				.b8(W2922D),
				.c(c2D209)
);

ninexnine_unit ninexnine_unit_4370(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2900E),
				.b1(W2901E),
				.b2(W2902E),
				.b3(W2910E),
				.b4(W2911E),
				.b5(W2912E),
				.b6(W2920E),
				.b7(W2921E),
				.b8(W2922E),
				.c(c2E209)
);

ninexnine_unit ninexnine_unit_4371(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2900F),
				.b1(W2901F),
				.b2(W2902F),
				.b3(W2910F),
				.b4(W2911F),
				.b5(W2912F),
				.b6(W2920F),
				.b7(W2921F),
				.b8(W2922F),
				.c(c2F209)
);

assign C2209=c20209+c21209+c22209+c23209+c24209+c25209+c26209+c27209+c28209+c29209+c2A209+c2B209+c2C209+c2D209+c2E209+c2F209;
assign A2209=(C2209>=0)?1:0;

assign P3209=A2209;

ninexnine_unit ninexnine_unit_4372(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20219)
);

ninexnine_unit ninexnine_unit_4373(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21219)
);

ninexnine_unit ninexnine_unit_4374(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22219)
);

ninexnine_unit ninexnine_unit_4375(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23219)
);

ninexnine_unit ninexnine_unit_4376(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24219)
);

ninexnine_unit ninexnine_unit_4377(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25219)
);

ninexnine_unit ninexnine_unit_4378(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26219)
);

ninexnine_unit ninexnine_unit_4379(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27219)
);

ninexnine_unit ninexnine_unit_4380(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W29008),
				.b1(W29018),
				.b2(W29028),
				.b3(W29108),
				.b4(W29118),
				.b5(W29128),
				.b6(W29208),
				.b7(W29218),
				.b8(W29228),
				.c(c28219)
);

ninexnine_unit ninexnine_unit_4381(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W29009),
				.b1(W29019),
				.b2(W29029),
				.b3(W29109),
				.b4(W29119),
				.b5(W29129),
				.b6(W29209),
				.b7(W29219),
				.b8(W29229),
				.c(c29219)
);

ninexnine_unit ninexnine_unit_4382(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2900A),
				.b1(W2901A),
				.b2(W2902A),
				.b3(W2910A),
				.b4(W2911A),
				.b5(W2912A),
				.b6(W2920A),
				.b7(W2921A),
				.b8(W2922A),
				.c(c2A219)
);

ninexnine_unit ninexnine_unit_4383(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2900B),
				.b1(W2901B),
				.b2(W2902B),
				.b3(W2910B),
				.b4(W2911B),
				.b5(W2912B),
				.b6(W2920B),
				.b7(W2921B),
				.b8(W2922B),
				.c(c2B219)
);

ninexnine_unit ninexnine_unit_4384(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2900C),
				.b1(W2901C),
				.b2(W2902C),
				.b3(W2910C),
				.b4(W2911C),
				.b5(W2912C),
				.b6(W2920C),
				.b7(W2921C),
				.b8(W2922C),
				.c(c2C219)
);

ninexnine_unit ninexnine_unit_4385(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2900D),
				.b1(W2901D),
				.b2(W2902D),
				.b3(W2910D),
				.b4(W2911D),
				.b5(W2912D),
				.b6(W2920D),
				.b7(W2921D),
				.b8(W2922D),
				.c(c2D219)
);

ninexnine_unit ninexnine_unit_4386(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2900E),
				.b1(W2901E),
				.b2(W2902E),
				.b3(W2910E),
				.b4(W2911E),
				.b5(W2912E),
				.b6(W2920E),
				.b7(W2921E),
				.b8(W2922E),
				.c(c2E219)
);

ninexnine_unit ninexnine_unit_4387(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2900F),
				.b1(W2901F),
				.b2(W2902F),
				.b3(W2910F),
				.b4(W2911F),
				.b5(W2912F),
				.b6(W2920F),
				.b7(W2921F),
				.b8(W2922F),
				.c(c2F219)
);

assign C2219=c20219+c21219+c22219+c23219+c24219+c25219+c26219+c27219+c28219+c29219+c2A219+c2B219+c2C219+c2D219+c2E219+c2F219;
assign A2219=(C2219>=0)?1:0;

assign P3219=A2219;

ninexnine_unit ninexnine_unit_4388(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W29000),
				.b1(W29010),
				.b2(W29020),
				.b3(W29100),
				.b4(W29110),
				.b5(W29120),
				.b6(W29200),
				.b7(W29210),
				.b8(W29220),
				.c(c20229)
);

ninexnine_unit ninexnine_unit_4389(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W29001),
				.b1(W29011),
				.b2(W29021),
				.b3(W29101),
				.b4(W29111),
				.b5(W29121),
				.b6(W29201),
				.b7(W29211),
				.b8(W29221),
				.c(c21229)
);

ninexnine_unit ninexnine_unit_4390(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W29002),
				.b1(W29012),
				.b2(W29022),
				.b3(W29102),
				.b4(W29112),
				.b5(W29122),
				.b6(W29202),
				.b7(W29212),
				.b8(W29222),
				.c(c22229)
);

ninexnine_unit ninexnine_unit_4391(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W29003),
				.b1(W29013),
				.b2(W29023),
				.b3(W29103),
				.b4(W29113),
				.b5(W29123),
				.b6(W29203),
				.b7(W29213),
				.b8(W29223),
				.c(c23229)
);

ninexnine_unit ninexnine_unit_4392(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W29004),
				.b1(W29014),
				.b2(W29024),
				.b3(W29104),
				.b4(W29114),
				.b5(W29124),
				.b6(W29204),
				.b7(W29214),
				.b8(W29224),
				.c(c24229)
);

ninexnine_unit ninexnine_unit_4393(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W29005),
				.b1(W29015),
				.b2(W29025),
				.b3(W29105),
				.b4(W29115),
				.b5(W29125),
				.b6(W29205),
				.b7(W29215),
				.b8(W29225),
				.c(c25229)
);

ninexnine_unit ninexnine_unit_4394(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W29006),
				.b1(W29016),
				.b2(W29026),
				.b3(W29106),
				.b4(W29116),
				.b5(W29126),
				.b6(W29206),
				.b7(W29216),
				.b8(W29226),
				.c(c26229)
);

ninexnine_unit ninexnine_unit_4395(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W29007),
				.b1(W29017),
				.b2(W29027),
				.b3(W29107),
				.b4(W29117),
				.b5(W29127),
				.b6(W29207),
				.b7(W29217),
				.b8(W29227),
				.c(c27229)
);

ninexnine_unit ninexnine_unit_4396(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W29008),
				.b1(W29018),
				.b2(W29028),
				.b3(W29108),
				.b4(W29118),
				.b5(W29128),
				.b6(W29208),
				.b7(W29218),
				.b8(W29228),
				.c(c28229)
);

ninexnine_unit ninexnine_unit_4397(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W29009),
				.b1(W29019),
				.b2(W29029),
				.b3(W29109),
				.b4(W29119),
				.b5(W29129),
				.b6(W29209),
				.b7(W29219),
				.b8(W29229),
				.c(c29229)
);

ninexnine_unit ninexnine_unit_4398(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2900A),
				.b1(W2901A),
				.b2(W2902A),
				.b3(W2910A),
				.b4(W2911A),
				.b5(W2912A),
				.b6(W2920A),
				.b7(W2921A),
				.b8(W2922A),
				.c(c2A229)
);

ninexnine_unit ninexnine_unit_4399(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2900B),
				.b1(W2901B),
				.b2(W2902B),
				.b3(W2910B),
				.b4(W2911B),
				.b5(W2912B),
				.b6(W2920B),
				.b7(W2921B),
				.b8(W2922B),
				.c(c2B229)
);

ninexnine_unit ninexnine_unit_4400(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2900C),
				.b1(W2901C),
				.b2(W2902C),
				.b3(W2910C),
				.b4(W2911C),
				.b5(W2912C),
				.b6(W2920C),
				.b7(W2921C),
				.b8(W2922C),
				.c(c2C229)
);

ninexnine_unit ninexnine_unit_4401(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2900D),
				.b1(W2901D),
				.b2(W2902D),
				.b3(W2910D),
				.b4(W2911D),
				.b5(W2912D),
				.b6(W2920D),
				.b7(W2921D),
				.b8(W2922D),
				.c(c2D229)
);

ninexnine_unit ninexnine_unit_4402(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2900E),
				.b1(W2901E),
				.b2(W2902E),
				.b3(W2910E),
				.b4(W2911E),
				.b5(W2912E),
				.b6(W2920E),
				.b7(W2921E),
				.b8(W2922E),
				.c(c2E229)
);

ninexnine_unit ninexnine_unit_4403(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2900F),
				.b1(W2901F),
				.b2(W2902F),
				.b3(W2910F),
				.b4(W2911F),
				.b5(W2912F),
				.b6(W2920F),
				.b7(W2921F),
				.b8(W2922F),
				.c(c2F229)
);

assign C2229=c20229+c21229+c22229+c23229+c24229+c25229+c26229+c27229+c28229+c29229+c2A229+c2B229+c2C229+c2D229+c2E229+c2F229;
assign A2229=(C2229>=0)?1:0;

assign P3229=A2229;

ninexnine_unit ninexnine_unit_4404(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2000A)
);

ninexnine_unit ninexnine_unit_4405(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2100A)
);

ninexnine_unit ninexnine_unit_4406(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2200A)
);

ninexnine_unit ninexnine_unit_4407(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2300A)
);

ninexnine_unit ninexnine_unit_4408(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2400A)
);

ninexnine_unit ninexnine_unit_4409(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2500A)
);

ninexnine_unit ninexnine_unit_4410(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2600A)
);

ninexnine_unit ninexnine_unit_4411(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2700A)
);

ninexnine_unit ninexnine_unit_4412(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2A008),
				.b1(W2A018),
				.b2(W2A028),
				.b3(W2A108),
				.b4(W2A118),
				.b5(W2A128),
				.b6(W2A208),
				.b7(W2A218),
				.b8(W2A228),
				.c(c2800A)
);

ninexnine_unit ninexnine_unit_4413(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2A009),
				.b1(W2A019),
				.b2(W2A029),
				.b3(W2A109),
				.b4(W2A119),
				.b5(W2A129),
				.b6(W2A209),
				.b7(W2A219),
				.b8(W2A229),
				.c(c2900A)
);

ninexnine_unit ninexnine_unit_4414(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2A00A),
				.b1(W2A01A),
				.b2(W2A02A),
				.b3(W2A10A),
				.b4(W2A11A),
				.b5(W2A12A),
				.b6(W2A20A),
				.b7(W2A21A),
				.b8(W2A22A),
				.c(c2A00A)
);

ninexnine_unit ninexnine_unit_4415(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2A00B),
				.b1(W2A01B),
				.b2(W2A02B),
				.b3(W2A10B),
				.b4(W2A11B),
				.b5(W2A12B),
				.b6(W2A20B),
				.b7(W2A21B),
				.b8(W2A22B),
				.c(c2B00A)
);

ninexnine_unit ninexnine_unit_4416(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2A00C),
				.b1(W2A01C),
				.b2(W2A02C),
				.b3(W2A10C),
				.b4(W2A11C),
				.b5(W2A12C),
				.b6(W2A20C),
				.b7(W2A21C),
				.b8(W2A22C),
				.c(c2C00A)
);

ninexnine_unit ninexnine_unit_4417(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2A00D),
				.b1(W2A01D),
				.b2(W2A02D),
				.b3(W2A10D),
				.b4(W2A11D),
				.b5(W2A12D),
				.b6(W2A20D),
				.b7(W2A21D),
				.b8(W2A22D),
				.c(c2D00A)
);

ninexnine_unit ninexnine_unit_4418(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2A00E),
				.b1(W2A01E),
				.b2(W2A02E),
				.b3(W2A10E),
				.b4(W2A11E),
				.b5(W2A12E),
				.b6(W2A20E),
				.b7(W2A21E),
				.b8(W2A22E),
				.c(c2E00A)
);

ninexnine_unit ninexnine_unit_4419(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2A00F),
				.b1(W2A01F),
				.b2(W2A02F),
				.b3(W2A10F),
				.b4(W2A11F),
				.b5(W2A12F),
				.b6(W2A20F),
				.b7(W2A21F),
				.b8(W2A22F),
				.c(c2F00A)
);

assign C200A=c2000A+c2100A+c2200A+c2300A+c2400A+c2500A+c2600A+c2700A+c2800A+c2900A+c2A00A+c2B00A+c2C00A+c2D00A+c2E00A+c2F00A;
assign A200A=(C200A>=0)?1:0;

assign P300A=A200A;

ninexnine_unit ninexnine_unit_4420(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2001A)
);

ninexnine_unit ninexnine_unit_4421(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2101A)
);

ninexnine_unit ninexnine_unit_4422(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2201A)
);

ninexnine_unit ninexnine_unit_4423(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2301A)
);

ninexnine_unit ninexnine_unit_4424(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2401A)
);

ninexnine_unit ninexnine_unit_4425(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2501A)
);

ninexnine_unit ninexnine_unit_4426(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2601A)
);

ninexnine_unit ninexnine_unit_4427(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2701A)
);

ninexnine_unit ninexnine_unit_4428(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2A008),
				.b1(W2A018),
				.b2(W2A028),
				.b3(W2A108),
				.b4(W2A118),
				.b5(W2A128),
				.b6(W2A208),
				.b7(W2A218),
				.b8(W2A228),
				.c(c2801A)
);

ninexnine_unit ninexnine_unit_4429(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2A009),
				.b1(W2A019),
				.b2(W2A029),
				.b3(W2A109),
				.b4(W2A119),
				.b5(W2A129),
				.b6(W2A209),
				.b7(W2A219),
				.b8(W2A229),
				.c(c2901A)
);

ninexnine_unit ninexnine_unit_4430(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2A00A),
				.b1(W2A01A),
				.b2(W2A02A),
				.b3(W2A10A),
				.b4(W2A11A),
				.b5(W2A12A),
				.b6(W2A20A),
				.b7(W2A21A),
				.b8(W2A22A),
				.c(c2A01A)
);

ninexnine_unit ninexnine_unit_4431(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2A00B),
				.b1(W2A01B),
				.b2(W2A02B),
				.b3(W2A10B),
				.b4(W2A11B),
				.b5(W2A12B),
				.b6(W2A20B),
				.b7(W2A21B),
				.b8(W2A22B),
				.c(c2B01A)
);

ninexnine_unit ninexnine_unit_4432(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2A00C),
				.b1(W2A01C),
				.b2(W2A02C),
				.b3(W2A10C),
				.b4(W2A11C),
				.b5(W2A12C),
				.b6(W2A20C),
				.b7(W2A21C),
				.b8(W2A22C),
				.c(c2C01A)
);

ninexnine_unit ninexnine_unit_4433(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2A00D),
				.b1(W2A01D),
				.b2(W2A02D),
				.b3(W2A10D),
				.b4(W2A11D),
				.b5(W2A12D),
				.b6(W2A20D),
				.b7(W2A21D),
				.b8(W2A22D),
				.c(c2D01A)
);

ninexnine_unit ninexnine_unit_4434(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2A00E),
				.b1(W2A01E),
				.b2(W2A02E),
				.b3(W2A10E),
				.b4(W2A11E),
				.b5(W2A12E),
				.b6(W2A20E),
				.b7(W2A21E),
				.b8(W2A22E),
				.c(c2E01A)
);

ninexnine_unit ninexnine_unit_4435(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2A00F),
				.b1(W2A01F),
				.b2(W2A02F),
				.b3(W2A10F),
				.b4(W2A11F),
				.b5(W2A12F),
				.b6(W2A20F),
				.b7(W2A21F),
				.b8(W2A22F),
				.c(c2F01A)
);

assign C201A=c2001A+c2101A+c2201A+c2301A+c2401A+c2501A+c2601A+c2701A+c2801A+c2901A+c2A01A+c2B01A+c2C01A+c2D01A+c2E01A+c2F01A;
assign A201A=(C201A>=0)?1:0;

assign P301A=A201A;

ninexnine_unit ninexnine_unit_4436(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2002A)
);

ninexnine_unit ninexnine_unit_4437(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2102A)
);

ninexnine_unit ninexnine_unit_4438(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2202A)
);

ninexnine_unit ninexnine_unit_4439(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2302A)
);

ninexnine_unit ninexnine_unit_4440(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2402A)
);

ninexnine_unit ninexnine_unit_4441(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2502A)
);

ninexnine_unit ninexnine_unit_4442(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2602A)
);

ninexnine_unit ninexnine_unit_4443(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2702A)
);

ninexnine_unit ninexnine_unit_4444(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2A008),
				.b1(W2A018),
				.b2(W2A028),
				.b3(W2A108),
				.b4(W2A118),
				.b5(W2A128),
				.b6(W2A208),
				.b7(W2A218),
				.b8(W2A228),
				.c(c2802A)
);

ninexnine_unit ninexnine_unit_4445(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2A009),
				.b1(W2A019),
				.b2(W2A029),
				.b3(W2A109),
				.b4(W2A119),
				.b5(W2A129),
				.b6(W2A209),
				.b7(W2A219),
				.b8(W2A229),
				.c(c2902A)
);

ninexnine_unit ninexnine_unit_4446(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2A00A),
				.b1(W2A01A),
				.b2(W2A02A),
				.b3(W2A10A),
				.b4(W2A11A),
				.b5(W2A12A),
				.b6(W2A20A),
				.b7(W2A21A),
				.b8(W2A22A),
				.c(c2A02A)
);

ninexnine_unit ninexnine_unit_4447(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2A00B),
				.b1(W2A01B),
				.b2(W2A02B),
				.b3(W2A10B),
				.b4(W2A11B),
				.b5(W2A12B),
				.b6(W2A20B),
				.b7(W2A21B),
				.b8(W2A22B),
				.c(c2B02A)
);

ninexnine_unit ninexnine_unit_4448(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2A00C),
				.b1(W2A01C),
				.b2(W2A02C),
				.b3(W2A10C),
				.b4(W2A11C),
				.b5(W2A12C),
				.b6(W2A20C),
				.b7(W2A21C),
				.b8(W2A22C),
				.c(c2C02A)
);

ninexnine_unit ninexnine_unit_4449(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2A00D),
				.b1(W2A01D),
				.b2(W2A02D),
				.b3(W2A10D),
				.b4(W2A11D),
				.b5(W2A12D),
				.b6(W2A20D),
				.b7(W2A21D),
				.b8(W2A22D),
				.c(c2D02A)
);

ninexnine_unit ninexnine_unit_4450(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2A00E),
				.b1(W2A01E),
				.b2(W2A02E),
				.b3(W2A10E),
				.b4(W2A11E),
				.b5(W2A12E),
				.b6(W2A20E),
				.b7(W2A21E),
				.b8(W2A22E),
				.c(c2E02A)
);

ninexnine_unit ninexnine_unit_4451(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2A00F),
				.b1(W2A01F),
				.b2(W2A02F),
				.b3(W2A10F),
				.b4(W2A11F),
				.b5(W2A12F),
				.b6(W2A20F),
				.b7(W2A21F),
				.b8(W2A22F),
				.c(c2F02A)
);

assign C202A=c2002A+c2102A+c2202A+c2302A+c2402A+c2502A+c2602A+c2702A+c2802A+c2902A+c2A02A+c2B02A+c2C02A+c2D02A+c2E02A+c2F02A;
assign A202A=(C202A>=0)?1:0;

assign P302A=A202A;

ninexnine_unit ninexnine_unit_4452(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2010A)
);

ninexnine_unit ninexnine_unit_4453(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2110A)
);

ninexnine_unit ninexnine_unit_4454(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2210A)
);

ninexnine_unit ninexnine_unit_4455(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2310A)
);

ninexnine_unit ninexnine_unit_4456(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2410A)
);

ninexnine_unit ninexnine_unit_4457(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2510A)
);

ninexnine_unit ninexnine_unit_4458(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2610A)
);

ninexnine_unit ninexnine_unit_4459(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2710A)
);

ninexnine_unit ninexnine_unit_4460(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2A008),
				.b1(W2A018),
				.b2(W2A028),
				.b3(W2A108),
				.b4(W2A118),
				.b5(W2A128),
				.b6(W2A208),
				.b7(W2A218),
				.b8(W2A228),
				.c(c2810A)
);

ninexnine_unit ninexnine_unit_4461(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2A009),
				.b1(W2A019),
				.b2(W2A029),
				.b3(W2A109),
				.b4(W2A119),
				.b5(W2A129),
				.b6(W2A209),
				.b7(W2A219),
				.b8(W2A229),
				.c(c2910A)
);

ninexnine_unit ninexnine_unit_4462(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2A00A),
				.b1(W2A01A),
				.b2(W2A02A),
				.b3(W2A10A),
				.b4(W2A11A),
				.b5(W2A12A),
				.b6(W2A20A),
				.b7(W2A21A),
				.b8(W2A22A),
				.c(c2A10A)
);

ninexnine_unit ninexnine_unit_4463(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2A00B),
				.b1(W2A01B),
				.b2(W2A02B),
				.b3(W2A10B),
				.b4(W2A11B),
				.b5(W2A12B),
				.b6(W2A20B),
				.b7(W2A21B),
				.b8(W2A22B),
				.c(c2B10A)
);

ninexnine_unit ninexnine_unit_4464(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2A00C),
				.b1(W2A01C),
				.b2(W2A02C),
				.b3(W2A10C),
				.b4(W2A11C),
				.b5(W2A12C),
				.b6(W2A20C),
				.b7(W2A21C),
				.b8(W2A22C),
				.c(c2C10A)
);

ninexnine_unit ninexnine_unit_4465(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2A00D),
				.b1(W2A01D),
				.b2(W2A02D),
				.b3(W2A10D),
				.b4(W2A11D),
				.b5(W2A12D),
				.b6(W2A20D),
				.b7(W2A21D),
				.b8(W2A22D),
				.c(c2D10A)
);

ninexnine_unit ninexnine_unit_4466(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2A00E),
				.b1(W2A01E),
				.b2(W2A02E),
				.b3(W2A10E),
				.b4(W2A11E),
				.b5(W2A12E),
				.b6(W2A20E),
				.b7(W2A21E),
				.b8(W2A22E),
				.c(c2E10A)
);

ninexnine_unit ninexnine_unit_4467(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2A00F),
				.b1(W2A01F),
				.b2(W2A02F),
				.b3(W2A10F),
				.b4(W2A11F),
				.b5(W2A12F),
				.b6(W2A20F),
				.b7(W2A21F),
				.b8(W2A22F),
				.c(c2F10A)
);

assign C210A=c2010A+c2110A+c2210A+c2310A+c2410A+c2510A+c2610A+c2710A+c2810A+c2910A+c2A10A+c2B10A+c2C10A+c2D10A+c2E10A+c2F10A;
assign A210A=(C210A>=0)?1:0;

assign P310A=A210A;

ninexnine_unit ninexnine_unit_4468(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2011A)
);

ninexnine_unit ninexnine_unit_4469(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2111A)
);

ninexnine_unit ninexnine_unit_4470(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2211A)
);

ninexnine_unit ninexnine_unit_4471(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2311A)
);

ninexnine_unit ninexnine_unit_4472(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2411A)
);

ninexnine_unit ninexnine_unit_4473(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2511A)
);

ninexnine_unit ninexnine_unit_4474(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2611A)
);

ninexnine_unit ninexnine_unit_4475(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2711A)
);

ninexnine_unit ninexnine_unit_4476(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2A008),
				.b1(W2A018),
				.b2(W2A028),
				.b3(W2A108),
				.b4(W2A118),
				.b5(W2A128),
				.b6(W2A208),
				.b7(W2A218),
				.b8(W2A228),
				.c(c2811A)
);

ninexnine_unit ninexnine_unit_4477(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2A009),
				.b1(W2A019),
				.b2(W2A029),
				.b3(W2A109),
				.b4(W2A119),
				.b5(W2A129),
				.b6(W2A209),
				.b7(W2A219),
				.b8(W2A229),
				.c(c2911A)
);

ninexnine_unit ninexnine_unit_4478(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2A00A),
				.b1(W2A01A),
				.b2(W2A02A),
				.b3(W2A10A),
				.b4(W2A11A),
				.b5(W2A12A),
				.b6(W2A20A),
				.b7(W2A21A),
				.b8(W2A22A),
				.c(c2A11A)
);

ninexnine_unit ninexnine_unit_4479(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2A00B),
				.b1(W2A01B),
				.b2(W2A02B),
				.b3(W2A10B),
				.b4(W2A11B),
				.b5(W2A12B),
				.b6(W2A20B),
				.b7(W2A21B),
				.b8(W2A22B),
				.c(c2B11A)
);

ninexnine_unit ninexnine_unit_4480(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2A00C),
				.b1(W2A01C),
				.b2(W2A02C),
				.b3(W2A10C),
				.b4(W2A11C),
				.b5(W2A12C),
				.b6(W2A20C),
				.b7(W2A21C),
				.b8(W2A22C),
				.c(c2C11A)
);

ninexnine_unit ninexnine_unit_4481(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2A00D),
				.b1(W2A01D),
				.b2(W2A02D),
				.b3(W2A10D),
				.b4(W2A11D),
				.b5(W2A12D),
				.b6(W2A20D),
				.b7(W2A21D),
				.b8(W2A22D),
				.c(c2D11A)
);

ninexnine_unit ninexnine_unit_4482(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2A00E),
				.b1(W2A01E),
				.b2(W2A02E),
				.b3(W2A10E),
				.b4(W2A11E),
				.b5(W2A12E),
				.b6(W2A20E),
				.b7(W2A21E),
				.b8(W2A22E),
				.c(c2E11A)
);

ninexnine_unit ninexnine_unit_4483(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2A00F),
				.b1(W2A01F),
				.b2(W2A02F),
				.b3(W2A10F),
				.b4(W2A11F),
				.b5(W2A12F),
				.b6(W2A20F),
				.b7(W2A21F),
				.b8(W2A22F),
				.c(c2F11A)
);

assign C211A=c2011A+c2111A+c2211A+c2311A+c2411A+c2511A+c2611A+c2711A+c2811A+c2911A+c2A11A+c2B11A+c2C11A+c2D11A+c2E11A+c2F11A;
assign A211A=(C211A>=0)?1:0;

assign P311A=A211A;

ninexnine_unit ninexnine_unit_4484(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2012A)
);

ninexnine_unit ninexnine_unit_4485(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2112A)
);

ninexnine_unit ninexnine_unit_4486(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2212A)
);

ninexnine_unit ninexnine_unit_4487(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2312A)
);

ninexnine_unit ninexnine_unit_4488(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2412A)
);

ninexnine_unit ninexnine_unit_4489(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2512A)
);

ninexnine_unit ninexnine_unit_4490(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2612A)
);

ninexnine_unit ninexnine_unit_4491(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2712A)
);

ninexnine_unit ninexnine_unit_4492(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2A008),
				.b1(W2A018),
				.b2(W2A028),
				.b3(W2A108),
				.b4(W2A118),
				.b5(W2A128),
				.b6(W2A208),
				.b7(W2A218),
				.b8(W2A228),
				.c(c2812A)
);

ninexnine_unit ninexnine_unit_4493(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2A009),
				.b1(W2A019),
				.b2(W2A029),
				.b3(W2A109),
				.b4(W2A119),
				.b5(W2A129),
				.b6(W2A209),
				.b7(W2A219),
				.b8(W2A229),
				.c(c2912A)
);

ninexnine_unit ninexnine_unit_4494(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2A00A),
				.b1(W2A01A),
				.b2(W2A02A),
				.b3(W2A10A),
				.b4(W2A11A),
				.b5(W2A12A),
				.b6(W2A20A),
				.b7(W2A21A),
				.b8(W2A22A),
				.c(c2A12A)
);

ninexnine_unit ninexnine_unit_4495(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2A00B),
				.b1(W2A01B),
				.b2(W2A02B),
				.b3(W2A10B),
				.b4(W2A11B),
				.b5(W2A12B),
				.b6(W2A20B),
				.b7(W2A21B),
				.b8(W2A22B),
				.c(c2B12A)
);

ninexnine_unit ninexnine_unit_4496(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2A00C),
				.b1(W2A01C),
				.b2(W2A02C),
				.b3(W2A10C),
				.b4(W2A11C),
				.b5(W2A12C),
				.b6(W2A20C),
				.b7(W2A21C),
				.b8(W2A22C),
				.c(c2C12A)
);

ninexnine_unit ninexnine_unit_4497(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2A00D),
				.b1(W2A01D),
				.b2(W2A02D),
				.b3(W2A10D),
				.b4(W2A11D),
				.b5(W2A12D),
				.b6(W2A20D),
				.b7(W2A21D),
				.b8(W2A22D),
				.c(c2D12A)
);

ninexnine_unit ninexnine_unit_4498(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2A00E),
				.b1(W2A01E),
				.b2(W2A02E),
				.b3(W2A10E),
				.b4(W2A11E),
				.b5(W2A12E),
				.b6(W2A20E),
				.b7(W2A21E),
				.b8(W2A22E),
				.c(c2E12A)
);

ninexnine_unit ninexnine_unit_4499(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2A00F),
				.b1(W2A01F),
				.b2(W2A02F),
				.b3(W2A10F),
				.b4(W2A11F),
				.b5(W2A12F),
				.b6(W2A20F),
				.b7(W2A21F),
				.b8(W2A22F),
				.c(c2F12A)
);

assign C212A=c2012A+c2112A+c2212A+c2312A+c2412A+c2512A+c2612A+c2712A+c2812A+c2912A+c2A12A+c2B12A+c2C12A+c2D12A+c2E12A+c2F12A;
assign A212A=(C212A>=0)?1:0;

assign P312A=A212A;

ninexnine_unit ninexnine_unit_4500(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2020A)
);

ninexnine_unit ninexnine_unit_4501(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2120A)
);

ninexnine_unit ninexnine_unit_4502(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2220A)
);

ninexnine_unit ninexnine_unit_4503(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2320A)
);

ninexnine_unit ninexnine_unit_4504(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2420A)
);

ninexnine_unit ninexnine_unit_4505(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2520A)
);

ninexnine_unit ninexnine_unit_4506(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2620A)
);

ninexnine_unit ninexnine_unit_4507(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2720A)
);

ninexnine_unit ninexnine_unit_4508(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2A008),
				.b1(W2A018),
				.b2(W2A028),
				.b3(W2A108),
				.b4(W2A118),
				.b5(W2A128),
				.b6(W2A208),
				.b7(W2A218),
				.b8(W2A228),
				.c(c2820A)
);

ninexnine_unit ninexnine_unit_4509(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2A009),
				.b1(W2A019),
				.b2(W2A029),
				.b3(W2A109),
				.b4(W2A119),
				.b5(W2A129),
				.b6(W2A209),
				.b7(W2A219),
				.b8(W2A229),
				.c(c2920A)
);

ninexnine_unit ninexnine_unit_4510(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2A00A),
				.b1(W2A01A),
				.b2(W2A02A),
				.b3(W2A10A),
				.b4(W2A11A),
				.b5(W2A12A),
				.b6(W2A20A),
				.b7(W2A21A),
				.b8(W2A22A),
				.c(c2A20A)
);

ninexnine_unit ninexnine_unit_4511(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2A00B),
				.b1(W2A01B),
				.b2(W2A02B),
				.b3(W2A10B),
				.b4(W2A11B),
				.b5(W2A12B),
				.b6(W2A20B),
				.b7(W2A21B),
				.b8(W2A22B),
				.c(c2B20A)
);

ninexnine_unit ninexnine_unit_4512(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2A00C),
				.b1(W2A01C),
				.b2(W2A02C),
				.b3(W2A10C),
				.b4(W2A11C),
				.b5(W2A12C),
				.b6(W2A20C),
				.b7(W2A21C),
				.b8(W2A22C),
				.c(c2C20A)
);

ninexnine_unit ninexnine_unit_4513(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2A00D),
				.b1(W2A01D),
				.b2(W2A02D),
				.b3(W2A10D),
				.b4(W2A11D),
				.b5(W2A12D),
				.b6(W2A20D),
				.b7(W2A21D),
				.b8(W2A22D),
				.c(c2D20A)
);

ninexnine_unit ninexnine_unit_4514(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2A00E),
				.b1(W2A01E),
				.b2(W2A02E),
				.b3(W2A10E),
				.b4(W2A11E),
				.b5(W2A12E),
				.b6(W2A20E),
				.b7(W2A21E),
				.b8(W2A22E),
				.c(c2E20A)
);

ninexnine_unit ninexnine_unit_4515(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2A00F),
				.b1(W2A01F),
				.b2(W2A02F),
				.b3(W2A10F),
				.b4(W2A11F),
				.b5(W2A12F),
				.b6(W2A20F),
				.b7(W2A21F),
				.b8(W2A22F),
				.c(c2F20A)
);

assign C220A=c2020A+c2120A+c2220A+c2320A+c2420A+c2520A+c2620A+c2720A+c2820A+c2920A+c2A20A+c2B20A+c2C20A+c2D20A+c2E20A+c2F20A;
assign A220A=(C220A>=0)?1:0;

assign P320A=A220A;

ninexnine_unit ninexnine_unit_4516(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2021A)
);

ninexnine_unit ninexnine_unit_4517(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2121A)
);

ninexnine_unit ninexnine_unit_4518(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2221A)
);

ninexnine_unit ninexnine_unit_4519(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2321A)
);

ninexnine_unit ninexnine_unit_4520(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2421A)
);

ninexnine_unit ninexnine_unit_4521(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2521A)
);

ninexnine_unit ninexnine_unit_4522(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2621A)
);

ninexnine_unit ninexnine_unit_4523(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2721A)
);

ninexnine_unit ninexnine_unit_4524(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2A008),
				.b1(W2A018),
				.b2(W2A028),
				.b3(W2A108),
				.b4(W2A118),
				.b5(W2A128),
				.b6(W2A208),
				.b7(W2A218),
				.b8(W2A228),
				.c(c2821A)
);

ninexnine_unit ninexnine_unit_4525(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2A009),
				.b1(W2A019),
				.b2(W2A029),
				.b3(W2A109),
				.b4(W2A119),
				.b5(W2A129),
				.b6(W2A209),
				.b7(W2A219),
				.b8(W2A229),
				.c(c2921A)
);

ninexnine_unit ninexnine_unit_4526(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2A00A),
				.b1(W2A01A),
				.b2(W2A02A),
				.b3(W2A10A),
				.b4(W2A11A),
				.b5(W2A12A),
				.b6(W2A20A),
				.b7(W2A21A),
				.b8(W2A22A),
				.c(c2A21A)
);

ninexnine_unit ninexnine_unit_4527(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2A00B),
				.b1(W2A01B),
				.b2(W2A02B),
				.b3(W2A10B),
				.b4(W2A11B),
				.b5(W2A12B),
				.b6(W2A20B),
				.b7(W2A21B),
				.b8(W2A22B),
				.c(c2B21A)
);

ninexnine_unit ninexnine_unit_4528(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2A00C),
				.b1(W2A01C),
				.b2(W2A02C),
				.b3(W2A10C),
				.b4(W2A11C),
				.b5(W2A12C),
				.b6(W2A20C),
				.b7(W2A21C),
				.b8(W2A22C),
				.c(c2C21A)
);

ninexnine_unit ninexnine_unit_4529(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2A00D),
				.b1(W2A01D),
				.b2(W2A02D),
				.b3(W2A10D),
				.b4(W2A11D),
				.b5(W2A12D),
				.b6(W2A20D),
				.b7(W2A21D),
				.b8(W2A22D),
				.c(c2D21A)
);

ninexnine_unit ninexnine_unit_4530(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2A00E),
				.b1(W2A01E),
				.b2(W2A02E),
				.b3(W2A10E),
				.b4(W2A11E),
				.b5(W2A12E),
				.b6(W2A20E),
				.b7(W2A21E),
				.b8(W2A22E),
				.c(c2E21A)
);

ninexnine_unit ninexnine_unit_4531(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2A00F),
				.b1(W2A01F),
				.b2(W2A02F),
				.b3(W2A10F),
				.b4(W2A11F),
				.b5(W2A12F),
				.b6(W2A20F),
				.b7(W2A21F),
				.b8(W2A22F),
				.c(c2F21A)
);

assign C221A=c2021A+c2121A+c2221A+c2321A+c2421A+c2521A+c2621A+c2721A+c2821A+c2921A+c2A21A+c2B21A+c2C21A+c2D21A+c2E21A+c2F21A;
assign A221A=(C221A>=0)?1:0;

assign P321A=A221A;

ninexnine_unit ninexnine_unit_4532(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2A000),
				.b1(W2A010),
				.b2(W2A020),
				.b3(W2A100),
				.b4(W2A110),
				.b5(W2A120),
				.b6(W2A200),
				.b7(W2A210),
				.b8(W2A220),
				.c(c2022A)
);

ninexnine_unit ninexnine_unit_4533(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2A001),
				.b1(W2A011),
				.b2(W2A021),
				.b3(W2A101),
				.b4(W2A111),
				.b5(W2A121),
				.b6(W2A201),
				.b7(W2A211),
				.b8(W2A221),
				.c(c2122A)
);

ninexnine_unit ninexnine_unit_4534(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2A002),
				.b1(W2A012),
				.b2(W2A022),
				.b3(W2A102),
				.b4(W2A112),
				.b5(W2A122),
				.b6(W2A202),
				.b7(W2A212),
				.b8(W2A222),
				.c(c2222A)
);

ninexnine_unit ninexnine_unit_4535(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2A003),
				.b1(W2A013),
				.b2(W2A023),
				.b3(W2A103),
				.b4(W2A113),
				.b5(W2A123),
				.b6(W2A203),
				.b7(W2A213),
				.b8(W2A223),
				.c(c2322A)
);

ninexnine_unit ninexnine_unit_4536(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2A004),
				.b1(W2A014),
				.b2(W2A024),
				.b3(W2A104),
				.b4(W2A114),
				.b5(W2A124),
				.b6(W2A204),
				.b7(W2A214),
				.b8(W2A224),
				.c(c2422A)
);

ninexnine_unit ninexnine_unit_4537(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2A005),
				.b1(W2A015),
				.b2(W2A025),
				.b3(W2A105),
				.b4(W2A115),
				.b5(W2A125),
				.b6(W2A205),
				.b7(W2A215),
				.b8(W2A225),
				.c(c2522A)
);

ninexnine_unit ninexnine_unit_4538(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2A006),
				.b1(W2A016),
				.b2(W2A026),
				.b3(W2A106),
				.b4(W2A116),
				.b5(W2A126),
				.b6(W2A206),
				.b7(W2A216),
				.b8(W2A226),
				.c(c2622A)
);

ninexnine_unit ninexnine_unit_4539(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2A007),
				.b1(W2A017),
				.b2(W2A027),
				.b3(W2A107),
				.b4(W2A117),
				.b5(W2A127),
				.b6(W2A207),
				.b7(W2A217),
				.b8(W2A227),
				.c(c2722A)
);

ninexnine_unit ninexnine_unit_4540(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2A008),
				.b1(W2A018),
				.b2(W2A028),
				.b3(W2A108),
				.b4(W2A118),
				.b5(W2A128),
				.b6(W2A208),
				.b7(W2A218),
				.b8(W2A228),
				.c(c2822A)
);

ninexnine_unit ninexnine_unit_4541(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2A009),
				.b1(W2A019),
				.b2(W2A029),
				.b3(W2A109),
				.b4(W2A119),
				.b5(W2A129),
				.b6(W2A209),
				.b7(W2A219),
				.b8(W2A229),
				.c(c2922A)
);

ninexnine_unit ninexnine_unit_4542(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2A00A),
				.b1(W2A01A),
				.b2(W2A02A),
				.b3(W2A10A),
				.b4(W2A11A),
				.b5(W2A12A),
				.b6(W2A20A),
				.b7(W2A21A),
				.b8(W2A22A),
				.c(c2A22A)
);

ninexnine_unit ninexnine_unit_4543(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2A00B),
				.b1(W2A01B),
				.b2(W2A02B),
				.b3(W2A10B),
				.b4(W2A11B),
				.b5(W2A12B),
				.b6(W2A20B),
				.b7(W2A21B),
				.b8(W2A22B),
				.c(c2B22A)
);

ninexnine_unit ninexnine_unit_4544(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2A00C),
				.b1(W2A01C),
				.b2(W2A02C),
				.b3(W2A10C),
				.b4(W2A11C),
				.b5(W2A12C),
				.b6(W2A20C),
				.b7(W2A21C),
				.b8(W2A22C),
				.c(c2C22A)
);

ninexnine_unit ninexnine_unit_4545(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2A00D),
				.b1(W2A01D),
				.b2(W2A02D),
				.b3(W2A10D),
				.b4(W2A11D),
				.b5(W2A12D),
				.b6(W2A20D),
				.b7(W2A21D),
				.b8(W2A22D),
				.c(c2D22A)
);

ninexnine_unit ninexnine_unit_4546(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2A00E),
				.b1(W2A01E),
				.b2(W2A02E),
				.b3(W2A10E),
				.b4(W2A11E),
				.b5(W2A12E),
				.b6(W2A20E),
				.b7(W2A21E),
				.b8(W2A22E),
				.c(c2E22A)
);

ninexnine_unit ninexnine_unit_4547(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2A00F),
				.b1(W2A01F),
				.b2(W2A02F),
				.b3(W2A10F),
				.b4(W2A11F),
				.b5(W2A12F),
				.b6(W2A20F),
				.b7(W2A21F),
				.b8(W2A22F),
				.c(c2F22A)
);

assign C222A=c2022A+c2122A+c2222A+c2322A+c2422A+c2522A+c2622A+c2722A+c2822A+c2922A+c2A22A+c2B22A+c2C22A+c2D22A+c2E22A+c2F22A;
assign A222A=(C222A>=0)?1:0;

assign P322A=A222A;

ninexnine_unit ninexnine_unit_4548(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2000B)
);

ninexnine_unit ninexnine_unit_4549(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2100B)
);

ninexnine_unit ninexnine_unit_4550(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2200B)
);

ninexnine_unit ninexnine_unit_4551(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2300B)
);

ninexnine_unit ninexnine_unit_4552(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2400B)
);

ninexnine_unit ninexnine_unit_4553(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2500B)
);

ninexnine_unit ninexnine_unit_4554(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2600B)
);

ninexnine_unit ninexnine_unit_4555(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2700B)
);

ninexnine_unit ninexnine_unit_4556(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2B008),
				.b1(W2B018),
				.b2(W2B028),
				.b3(W2B108),
				.b4(W2B118),
				.b5(W2B128),
				.b6(W2B208),
				.b7(W2B218),
				.b8(W2B228),
				.c(c2800B)
);

ninexnine_unit ninexnine_unit_4557(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2B009),
				.b1(W2B019),
				.b2(W2B029),
				.b3(W2B109),
				.b4(W2B119),
				.b5(W2B129),
				.b6(W2B209),
				.b7(W2B219),
				.b8(W2B229),
				.c(c2900B)
);

ninexnine_unit ninexnine_unit_4558(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2B00A),
				.b1(W2B01A),
				.b2(W2B02A),
				.b3(W2B10A),
				.b4(W2B11A),
				.b5(W2B12A),
				.b6(W2B20A),
				.b7(W2B21A),
				.b8(W2B22A),
				.c(c2A00B)
);

ninexnine_unit ninexnine_unit_4559(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2B00B),
				.b1(W2B01B),
				.b2(W2B02B),
				.b3(W2B10B),
				.b4(W2B11B),
				.b5(W2B12B),
				.b6(W2B20B),
				.b7(W2B21B),
				.b8(W2B22B),
				.c(c2B00B)
);

ninexnine_unit ninexnine_unit_4560(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2B00C),
				.b1(W2B01C),
				.b2(W2B02C),
				.b3(W2B10C),
				.b4(W2B11C),
				.b5(W2B12C),
				.b6(W2B20C),
				.b7(W2B21C),
				.b8(W2B22C),
				.c(c2C00B)
);

ninexnine_unit ninexnine_unit_4561(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2B00D),
				.b1(W2B01D),
				.b2(W2B02D),
				.b3(W2B10D),
				.b4(W2B11D),
				.b5(W2B12D),
				.b6(W2B20D),
				.b7(W2B21D),
				.b8(W2B22D),
				.c(c2D00B)
);

ninexnine_unit ninexnine_unit_4562(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2B00E),
				.b1(W2B01E),
				.b2(W2B02E),
				.b3(W2B10E),
				.b4(W2B11E),
				.b5(W2B12E),
				.b6(W2B20E),
				.b7(W2B21E),
				.b8(W2B22E),
				.c(c2E00B)
);

ninexnine_unit ninexnine_unit_4563(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2B00F),
				.b1(W2B01F),
				.b2(W2B02F),
				.b3(W2B10F),
				.b4(W2B11F),
				.b5(W2B12F),
				.b6(W2B20F),
				.b7(W2B21F),
				.b8(W2B22F),
				.c(c2F00B)
);

assign C200B=c2000B+c2100B+c2200B+c2300B+c2400B+c2500B+c2600B+c2700B+c2800B+c2900B+c2A00B+c2B00B+c2C00B+c2D00B+c2E00B+c2F00B;
assign A200B=(C200B>=0)?1:0;

assign P300B=A200B;

ninexnine_unit ninexnine_unit_4564(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2001B)
);

ninexnine_unit ninexnine_unit_4565(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2101B)
);

ninexnine_unit ninexnine_unit_4566(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2201B)
);

ninexnine_unit ninexnine_unit_4567(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2301B)
);

ninexnine_unit ninexnine_unit_4568(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2401B)
);

ninexnine_unit ninexnine_unit_4569(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2501B)
);

ninexnine_unit ninexnine_unit_4570(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2601B)
);

ninexnine_unit ninexnine_unit_4571(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2701B)
);

ninexnine_unit ninexnine_unit_4572(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2B008),
				.b1(W2B018),
				.b2(W2B028),
				.b3(W2B108),
				.b4(W2B118),
				.b5(W2B128),
				.b6(W2B208),
				.b7(W2B218),
				.b8(W2B228),
				.c(c2801B)
);

ninexnine_unit ninexnine_unit_4573(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2B009),
				.b1(W2B019),
				.b2(W2B029),
				.b3(W2B109),
				.b4(W2B119),
				.b5(W2B129),
				.b6(W2B209),
				.b7(W2B219),
				.b8(W2B229),
				.c(c2901B)
);

ninexnine_unit ninexnine_unit_4574(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2B00A),
				.b1(W2B01A),
				.b2(W2B02A),
				.b3(W2B10A),
				.b4(W2B11A),
				.b5(W2B12A),
				.b6(W2B20A),
				.b7(W2B21A),
				.b8(W2B22A),
				.c(c2A01B)
);

ninexnine_unit ninexnine_unit_4575(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2B00B),
				.b1(W2B01B),
				.b2(W2B02B),
				.b3(W2B10B),
				.b4(W2B11B),
				.b5(W2B12B),
				.b6(W2B20B),
				.b7(W2B21B),
				.b8(W2B22B),
				.c(c2B01B)
);

ninexnine_unit ninexnine_unit_4576(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2B00C),
				.b1(W2B01C),
				.b2(W2B02C),
				.b3(W2B10C),
				.b4(W2B11C),
				.b5(W2B12C),
				.b6(W2B20C),
				.b7(W2B21C),
				.b8(W2B22C),
				.c(c2C01B)
);

ninexnine_unit ninexnine_unit_4577(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2B00D),
				.b1(W2B01D),
				.b2(W2B02D),
				.b3(W2B10D),
				.b4(W2B11D),
				.b5(W2B12D),
				.b6(W2B20D),
				.b7(W2B21D),
				.b8(W2B22D),
				.c(c2D01B)
);

ninexnine_unit ninexnine_unit_4578(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2B00E),
				.b1(W2B01E),
				.b2(W2B02E),
				.b3(W2B10E),
				.b4(W2B11E),
				.b5(W2B12E),
				.b6(W2B20E),
				.b7(W2B21E),
				.b8(W2B22E),
				.c(c2E01B)
);

ninexnine_unit ninexnine_unit_4579(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2B00F),
				.b1(W2B01F),
				.b2(W2B02F),
				.b3(W2B10F),
				.b4(W2B11F),
				.b5(W2B12F),
				.b6(W2B20F),
				.b7(W2B21F),
				.b8(W2B22F),
				.c(c2F01B)
);

assign C201B=c2001B+c2101B+c2201B+c2301B+c2401B+c2501B+c2601B+c2701B+c2801B+c2901B+c2A01B+c2B01B+c2C01B+c2D01B+c2E01B+c2F01B;
assign A201B=(C201B>=0)?1:0;

assign P301B=A201B;

ninexnine_unit ninexnine_unit_4580(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2002B)
);

ninexnine_unit ninexnine_unit_4581(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2102B)
);

ninexnine_unit ninexnine_unit_4582(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2202B)
);

ninexnine_unit ninexnine_unit_4583(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2302B)
);

ninexnine_unit ninexnine_unit_4584(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2402B)
);

ninexnine_unit ninexnine_unit_4585(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2502B)
);

ninexnine_unit ninexnine_unit_4586(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2602B)
);

ninexnine_unit ninexnine_unit_4587(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2702B)
);

ninexnine_unit ninexnine_unit_4588(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2B008),
				.b1(W2B018),
				.b2(W2B028),
				.b3(W2B108),
				.b4(W2B118),
				.b5(W2B128),
				.b6(W2B208),
				.b7(W2B218),
				.b8(W2B228),
				.c(c2802B)
);

ninexnine_unit ninexnine_unit_4589(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2B009),
				.b1(W2B019),
				.b2(W2B029),
				.b3(W2B109),
				.b4(W2B119),
				.b5(W2B129),
				.b6(W2B209),
				.b7(W2B219),
				.b8(W2B229),
				.c(c2902B)
);

ninexnine_unit ninexnine_unit_4590(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2B00A),
				.b1(W2B01A),
				.b2(W2B02A),
				.b3(W2B10A),
				.b4(W2B11A),
				.b5(W2B12A),
				.b6(W2B20A),
				.b7(W2B21A),
				.b8(W2B22A),
				.c(c2A02B)
);

ninexnine_unit ninexnine_unit_4591(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2B00B),
				.b1(W2B01B),
				.b2(W2B02B),
				.b3(W2B10B),
				.b4(W2B11B),
				.b5(W2B12B),
				.b6(W2B20B),
				.b7(W2B21B),
				.b8(W2B22B),
				.c(c2B02B)
);

ninexnine_unit ninexnine_unit_4592(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2B00C),
				.b1(W2B01C),
				.b2(W2B02C),
				.b3(W2B10C),
				.b4(W2B11C),
				.b5(W2B12C),
				.b6(W2B20C),
				.b7(W2B21C),
				.b8(W2B22C),
				.c(c2C02B)
);

ninexnine_unit ninexnine_unit_4593(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2B00D),
				.b1(W2B01D),
				.b2(W2B02D),
				.b3(W2B10D),
				.b4(W2B11D),
				.b5(W2B12D),
				.b6(W2B20D),
				.b7(W2B21D),
				.b8(W2B22D),
				.c(c2D02B)
);

ninexnine_unit ninexnine_unit_4594(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2B00E),
				.b1(W2B01E),
				.b2(W2B02E),
				.b3(W2B10E),
				.b4(W2B11E),
				.b5(W2B12E),
				.b6(W2B20E),
				.b7(W2B21E),
				.b8(W2B22E),
				.c(c2E02B)
);

ninexnine_unit ninexnine_unit_4595(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2B00F),
				.b1(W2B01F),
				.b2(W2B02F),
				.b3(W2B10F),
				.b4(W2B11F),
				.b5(W2B12F),
				.b6(W2B20F),
				.b7(W2B21F),
				.b8(W2B22F),
				.c(c2F02B)
);

assign C202B=c2002B+c2102B+c2202B+c2302B+c2402B+c2502B+c2602B+c2702B+c2802B+c2902B+c2A02B+c2B02B+c2C02B+c2D02B+c2E02B+c2F02B;
assign A202B=(C202B>=0)?1:0;

assign P302B=A202B;

ninexnine_unit ninexnine_unit_4596(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2010B)
);

ninexnine_unit ninexnine_unit_4597(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2110B)
);

ninexnine_unit ninexnine_unit_4598(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2210B)
);

ninexnine_unit ninexnine_unit_4599(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2310B)
);

ninexnine_unit ninexnine_unit_4600(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2410B)
);

ninexnine_unit ninexnine_unit_4601(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2510B)
);

ninexnine_unit ninexnine_unit_4602(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2610B)
);

ninexnine_unit ninexnine_unit_4603(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2710B)
);

ninexnine_unit ninexnine_unit_4604(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2B008),
				.b1(W2B018),
				.b2(W2B028),
				.b3(W2B108),
				.b4(W2B118),
				.b5(W2B128),
				.b6(W2B208),
				.b7(W2B218),
				.b8(W2B228),
				.c(c2810B)
);

ninexnine_unit ninexnine_unit_4605(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2B009),
				.b1(W2B019),
				.b2(W2B029),
				.b3(W2B109),
				.b4(W2B119),
				.b5(W2B129),
				.b6(W2B209),
				.b7(W2B219),
				.b8(W2B229),
				.c(c2910B)
);

ninexnine_unit ninexnine_unit_4606(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2B00A),
				.b1(W2B01A),
				.b2(W2B02A),
				.b3(W2B10A),
				.b4(W2B11A),
				.b5(W2B12A),
				.b6(W2B20A),
				.b7(W2B21A),
				.b8(W2B22A),
				.c(c2A10B)
);

ninexnine_unit ninexnine_unit_4607(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2B00B),
				.b1(W2B01B),
				.b2(W2B02B),
				.b3(W2B10B),
				.b4(W2B11B),
				.b5(W2B12B),
				.b6(W2B20B),
				.b7(W2B21B),
				.b8(W2B22B),
				.c(c2B10B)
);

ninexnine_unit ninexnine_unit_4608(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2B00C),
				.b1(W2B01C),
				.b2(W2B02C),
				.b3(W2B10C),
				.b4(W2B11C),
				.b5(W2B12C),
				.b6(W2B20C),
				.b7(W2B21C),
				.b8(W2B22C),
				.c(c2C10B)
);

ninexnine_unit ninexnine_unit_4609(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2B00D),
				.b1(W2B01D),
				.b2(W2B02D),
				.b3(W2B10D),
				.b4(W2B11D),
				.b5(W2B12D),
				.b6(W2B20D),
				.b7(W2B21D),
				.b8(W2B22D),
				.c(c2D10B)
);

ninexnine_unit ninexnine_unit_4610(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2B00E),
				.b1(W2B01E),
				.b2(W2B02E),
				.b3(W2B10E),
				.b4(W2B11E),
				.b5(W2B12E),
				.b6(W2B20E),
				.b7(W2B21E),
				.b8(W2B22E),
				.c(c2E10B)
);

ninexnine_unit ninexnine_unit_4611(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2B00F),
				.b1(W2B01F),
				.b2(W2B02F),
				.b3(W2B10F),
				.b4(W2B11F),
				.b5(W2B12F),
				.b6(W2B20F),
				.b7(W2B21F),
				.b8(W2B22F),
				.c(c2F10B)
);

assign C210B=c2010B+c2110B+c2210B+c2310B+c2410B+c2510B+c2610B+c2710B+c2810B+c2910B+c2A10B+c2B10B+c2C10B+c2D10B+c2E10B+c2F10B;
assign A210B=(C210B>=0)?1:0;

assign P310B=A210B;

ninexnine_unit ninexnine_unit_4612(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2011B)
);

ninexnine_unit ninexnine_unit_4613(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2111B)
);

ninexnine_unit ninexnine_unit_4614(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2211B)
);

ninexnine_unit ninexnine_unit_4615(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2311B)
);

ninexnine_unit ninexnine_unit_4616(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2411B)
);

ninexnine_unit ninexnine_unit_4617(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2511B)
);

ninexnine_unit ninexnine_unit_4618(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2611B)
);

ninexnine_unit ninexnine_unit_4619(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2711B)
);

ninexnine_unit ninexnine_unit_4620(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2B008),
				.b1(W2B018),
				.b2(W2B028),
				.b3(W2B108),
				.b4(W2B118),
				.b5(W2B128),
				.b6(W2B208),
				.b7(W2B218),
				.b8(W2B228),
				.c(c2811B)
);

ninexnine_unit ninexnine_unit_4621(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2B009),
				.b1(W2B019),
				.b2(W2B029),
				.b3(W2B109),
				.b4(W2B119),
				.b5(W2B129),
				.b6(W2B209),
				.b7(W2B219),
				.b8(W2B229),
				.c(c2911B)
);

ninexnine_unit ninexnine_unit_4622(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2B00A),
				.b1(W2B01A),
				.b2(W2B02A),
				.b3(W2B10A),
				.b4(W2B11A),
				.b5(W2B12A),
				.b6(W2B20A),
				.b7(W2B21A),
				.b8(W2B22A),
				.c(c2A11B)
);

ninexnine_unit ninexnine_unit_4623(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2B00B),
				.b1(W2B01B),
				.b2(W2B02B),
				.b3(W2B10B),
				.b4(W2B11B),
				.b5(W2B12B),
				.b6(W2B20B),
				.b7(W2B21B),
				.b8(W2B22B),
				.c(c2B11B)
);

ninexnine_unit ninexnine_unit_4624(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2B00C),
				.b1(W2B01C),
				.b2(W2B02C),
				.b3(W2B10C),
				.b4(W2B11C),
				.b5(W2B12C),
				.b6(W2B20C),
				.b7(W2B21C),
				.b8(W2B22C),
				.c(c2C11B)
);

ninexnine_unit ninexnine_unit_4625(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2B00D),
				.b1(W2B01D),
				.b2(W2B02D),
				.b3(W2B10D),
				.b4(W2B11D),
				.b5(W2B12D),
				.b6(W2B20D),
				.b7(W2B21D),
				.b8(W2B22D),
				.c(c2D11B)
);

ninexnine_unit ninexnine_unit_4626(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2B00E),
				.b1(W2B01E),
				.b2(W2B02E),
				.b3(W2B10E),
				.b4(W2B11E),
				.b5(W2B12E),
				.b6(W2B20E),
				.b7(W2B21E),
				.b8(W2B22E),
				.c(c2E11B)
);

ninexnine_unit ninexnine_unit_4627(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2B00F),
				.b1(W2B01F),
				.b2(W2B02F),
				.b3(W2B10F),
				.b4(W2B11F),
				.b5(W2B12F),
				.b6(W2B20F),
				.b7(W2B21F),
				.b8(W2B22F),
				.c(c2F11B)
);

assign C211B=c2011B+c2111B+c2211B+c2311B+c2411B+c2511B+c2611B+c2711B+c2811B+c2911B+c2A11B+c2B11B+c2C11B+c2D11B+c2E11B+c2F11B;
assign A211B=(C211B>=0)?1:0;

assign P311B=A211B;

ninexnine_unit ninexnine_unit_4628(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2012B)
);

ninexnine_unit ninexnine_unit_4629(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2112B)
);

ninexnine_unit ninexnine_unit_4630(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2212B)
);

ninexnine_unit ninexnine_unit_4631(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2312B)
);

ninexnine_unit ninexnine_unit_4632(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2412B)
);

ninexnine_unit ninexnine_unit_4633(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2512B)
);

ninexnine_unit ninexnine_unit_4634(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2612B)
);

ninexnine_unit ninexnine_unit_4635(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2712B)
);

ninexnine_unit ninexnine_unit_4636(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2B008),
				.b1(W2B018),
				.b2(W2B028),
				.b3(W2B108),
				.b4(W2B118),
				.b5(W2B128),
				.b6(W2B208),
				.b7(W2B218),
				.b8(W2B228),
				.c(c2812B)
);

ninexnine_unit ninexnine_unit_4637(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2B009),
				.b1(W2B019),
				.b2(W2B029),
				.b3(W2B109),
				.b4(W2B119),
				.b5(W2B129),
				.b6(W2B209),
				.b7(W2B219),
				.b8(W2B229),
				.c(c2912B)
);

ninexnine_unit ninexnine_unit_4638(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2B00A),
				.b1(W2B01A),
				.b2(W2B02A),
				.b3(W2B10A),
				.b4(W2B11A),
				.b5(W2B12A),
				.b6(W2B20A),
				.b7(W2B21A),
				.b8(W2B22A),
				.c(c2A12B)
);

ninexnine_unit ninexnine_unit_4639(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2B00B),
				.b1(W2B01B),
				.b2(W2B02B),
				.b3(W2B10B),
				.b4(W2B11B),
				.b5(W2B12B),
				.b6(W2B20B),
				.b7(W2B21B),
				.b8(W2B22B),
				.c(c2B12B)
);

ninexnine_unit ninexnine_unit_4640(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2B00C),
				.b1(W2B01C),
				.b2(W2B02C),
				.b3(W2B10C),
				.b4(W2B11C),
				.b5(W2B12C),
				.b6(W2B20C),
				.b7(W2B21C),
				.b8(W2B22C),
				.c(c2C12B)
);

ninexnine_unit ninexnine_unit_4641(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2B00D),
				.b1(W2B01D),
				.b2(W2B02D),
				.b3(W2B10D),
				.b4(W2B11D),
				.b5(W2B12D),
				.b6(W2B20D),
				.b7(W2B21D),
				.b8(W2B22D),
				.c(c2D12B)
);

ninexnine_unit ninexnine_unit_4642(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2B00E),
				.b1(W2B01E),
				.b2(W2B02E),
				.b3(W2B10E),
				.b4(W2B11E),
				.b5(W2B12E),
				.b6(W2B20E),
				.b7(W2B21E),
				.b8(W2B22E),
				.c(c2E12B)
);

ninexnine_unit ninexnine_unit_4643(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2B00F),
				.b1(W2B01F),
				.b2(W2B02F),
				.b3(W2B10F),
				.b4(W2B11F),
				.b5(W2B12F),
				.b6(W2B20F),
				.b7(W2B21F),
				.b8(W2B22F),
				.c(c2F12B)
);

assign C212B=c2012B+c2112B+c2212B+c2312B+c2412B+c2512B+c2612B+c2712B+c2812B+c2912B+c2A12B+c2B12B+c2C12B+c2D12B+c2E12B+c2F12B;
assign A212B=(C212B>=0)?1:0;

assign P312B=A212B;

ninexnine_unit ninexnine_unit_4644(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2020B)
);

ninexnine_unit ninexnine_unit_4645(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2120B)
);

ninexnine_unit ninexnine_unit_4646(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2220B)
);

ninexnine_unit ninexnine_unit_4647(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2320B)
);

ninexnine_unit ninexnine_unit_4648(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2420B)
);

ninexnine_unit ninexnine_unit_4649(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2520B)
);

ninexnine_unit ninexnine_unit_4650(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2620B)
);

ninexnine_unit ninexnine_unit_4651(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2720B)
);

ninexnine_unit ninexnine_unit_4652(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2B008),
				.b1(W2B018),
				.b2(W2B028),
				.b3(W2B108),
				.b4(W2B118),
				.b5(W2B128),
				.b6(W2B208),
				.b7(W2B218),
				.b8(W2B228),
				.c(c2820B)
);

ninexnine_unit ninexnine_unit_4653(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2B009),
				.b1(W2B019),
				.b2(W2B029),
				.b3(W2B109),
				.b4(W2B119),
				.b5(W2B129),
				.b6(W2B209),
				.b7(W2B219),
				.b8(W2B229),
				.c(c2920B)
);

ninexnine_unit ninexnine_unit_4654(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2B00A),
				.b1(W2B01A),
				.b2(W2B02A),
				.b3(W2B10A),
				.b4(W2B11A),
				.b5(W2B12A),
				.b6(W2B20A),
				.b7(W2B21A),
				.b8(W2B22A),
				.c(c2A20B)
);

ninexnine_unit ninexnine_unit_4655(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2B00B),
				.b1(W2B01B),
				.b2(W2B02B),
				.b3(W2B10B),
				.b4(W2B11B),
				.b5(W2B12B),
				.b6(W2B20B),
				.b7(W2B21B),
				.b8(W2B22B),
				.c(c2B20B)
);

ninexnine_unit ninexnine_unit_4656(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2B00C),
				.b1(W2B01C),
				.b2(W2B02C),
				.b3(W2B10C),
				.b4(W2B11C),
				.b5(W2B12C),
				.b6(W2B20C),
				.b7(W2B21C),
				.b8(W2B22C),
				.c(c2C20B)
);

ninexnine_unit ninexnine_unit_4657(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2B00D),
				.b1(W2B01D),
				.b2(W2B02D),
				.b3(W2B10D),
				.b4(W2B11D),
				.b5(W2B12D),
				.b6(W2B20D),
				.b7(W2B21D),
				.b8(W2B22D),
				.c(c2D20B)
);

ninexnine_unit ninexnine_unit_4658(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2B00E),
				.b1(W2B01E),
				.b2(W2B02E),
				.b3(W2B10E),
				.b4(W2B11E),
				.b5(W2B12E),
				.b6(W2B20E),
				.b7(W2B21E),
				.b8(W2B22E),
				.c(c2E20B)
);

ninexnine_unit ninexnine_unit_4659(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2B00F),
				.b1(W2B01F),
				.b2(W2B02F),
				.b3(W2B10F),
				.b4(W2B11F),
				.b5(W2B12F),
				.b6(W2B20F),
				.b7(W2B21F),
				.b8(W2B22F),
				.c(c2F20B)
);

assign C220B=c2020B+c2120B+c2220B+c2320B+c2420B+c2520B+c2620B+c2720B+c2820B+c2920B+c2A20B+c2B20B+c2C20B+c2D20B+c2E20B+c2F20B;
assign A220B=(C220B>=0)?1:0;

assign P320B=A220B;

ninexnine_unit ninexnine_unit_4660(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2021B)
);

ninexnine_unit ninexnine_unit_4661(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2121B)
);

ninexnine_unit ninexnine_unit_4662(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2221B)
);

ninexnine_unit ninexnine_unit_4663(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2321B)
);

ninexnine_unit ninexnine_unit_4664(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2421B)
);

ninexnine_unit ninexnine_unit_4665(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2521B)
);

ninexnine_unit ninexnine_unit_4666(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2621B)
);

ninexnine_unit ninexnine_unit_4667(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2721B)
);

ninexnine_unit ninexnine_unit_4668(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2B008),
				.b1(W2B018),
				.b2(W2B028),
				.b3(W2B108),
				.b4(W2B118),
				.b5(W2B128),
				.b6(W2B208),
				.b7(W2B218),
				.b8(W2B228),
				.c(c2821B)
);

ninexnine_unit ninexnine_unit_4669(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2B009),
				.b1(W2B019),
				.b2(W2B029),
				.b3(W2B109),
				.b4(W2B119),
				.b5(W2B129),
				.b6(W2B209),
				.b7(W2B219),
				.b8(W2B229),
				.c(c2921B)
);

ninexnine_unit ninexnine_unit_4670(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2B00A),
				.b1(W2B01A),
				.b2(W2B02A),
				.b3(W2B10A),
				.b4(W2B11A),
				.b5(W2B12A),
				.b6(W2B20A),
				.b7(W2B21A),
				.b8(W2B22A),
				.c(c2A21B)
);

ninexnine_unit ninexnine_unit_4671(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2B00B),
				.b1(W2B01B),
				.b2(W2B02B),
				.b3(W2B10B),
				.b4(W2B11B),
				.b5(W2B12B),
				.b6(W2B20B),
				.b7(W2B21B),
				.b8(W2B22B),
				.c(c2B21B)
);

ninexnine_unit ninexnine_unit_4672(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2B00C),
				.b1(W2B01C),
				.b2(W2B02C),
				.b3(W2B10C),
				.b4(W2B11C),
				.b5(W2B12C),
				.b6(W2B20C),
				.b7(W2B21C),
				.b8(W2B22C),
				.c(c2C21B)
);

ninexnine_unit ninexnine_unit_4673(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2B00D),
				.b1(W2B01D),
				.b2(W2B02D),
				.b3(W2B10D),
				.b4(W2B11D),
				.b5(W2B12D),
				.b6(W2B20D),
				.b7(W2B21D),
				.b8(W2B22D),
				.c(c2D21B)
);

ninexnine_unit ninexnine_unit_4674(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2B00E),
				.b1(W2B01E),
				.b2(W2B02E),
				.b3(W2B10E),
				.b4(W2B11E),
				.b5(W2B12E),
				.b6(W2B20E),
				.b7(W2B21E),
				.b8(W2B22E),
				.c(c2E21B)
);

ninexnine_unit ninexnine_unit_4675(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2B00F),
				.b1(W2B01F),
				.b2(W2B02F),
				.b3(W2B10F),
				.b4(W2B11F),
				.b5(W2B12F),
				.b6(W2B20F),
				.b7(W2B21F),
				.b8(W2B22F),
				.c(c2F21B)
);

assign C221B=c2021B+c2121B+c2221B+c2321B+c2421B+c2521B+c2621B+c2721B+c2821B+c2921B+c2A21B+c2B21B+c2C21B+c2D21B+c2E21B+c2F21B;
assign A221B=(C221B>=0)?1:0;

assign P321B=A221B;

ninexnine_unit ninexnine_unit_4676(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2B000),
				.b1(W2B010),
				.b2(W2B020),
				.b3(W2B100),
				.b4(W2B110),
				.b5(W2B120),
				.b6(W2B200),
				.b7(W2B210),
				.b8(W2B220),
				.c(c2022B)
);

ninexnine_unit ninexnine_unit_4677(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2B001),
				.b1(W2B011),
				.b2(W2B021),
				.b3(W2B101),
				.b4(W2B111),
				.b5(W2B121),
				.b6(W2B201),
				.b7(W2B211),
				.b8(W2B221),
				.c(c2122B)
);

ninexnine_unit ninexnine_unit_4678(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2B002),
				.b1(W2B012),
				.b2(W2B022),
				.b3(W2B102),
				.b4(W2B112),
				.b5(W2B122),
				.b6(W2B202),
				.b7(W2B212),
				.b8(W2B222),
				.c(c2222B)
);

ninexnine_unit ninexnine_unit_4679(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2B003),
				.b1(W2B013),
				.b2(W2B023),
				.b3(W2B103),
				.b4(W2B113),
				.b5(W2B123),
				.b6(W2B203),
				.b7(W2B213),
				.b8(W2B223),
				.c(c2322B)
);

ninexnine_unit ninexnine_unit_4680(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2B004),
				.b1(W2B014),
				.b2(W2B024),
				.b3(W2B104),
				.b4(W2B114),
				.b5(W2B124),
				.b6(W2B204),
				.b7(W2B214),
				.b8(W2B224),
				.c(c2422B)
);

ninexnine_unit ninexnine_unit_4681(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2B005),
				.b1(W2B015),
				.b2(W2B025),
				.b3(W2B105),
				.b4(W2B115),
				.b5(W2B125),
				.b6(W2B205),
				.b7(W2B215),
				.b8(W2B225),
				.c(c2522B)
);

ninexnine_unit ninexnine_unit_4682(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2B006),
				.b1(W2B016),
				.b2(W2B026),
				.b3(W2B106),
				.b4(W2B116),
				.b5(W2B126),
				.b6(W2B206),
				.b7(W2B216),
				.b8(W2B226),
				.c(c2622B)
);

ninexnine_unit ninexnine_unit_4683(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2B007),
				.b1(W2B017),
				.b2(W2B027),
				.b3(W2B107),
				.b4(W2B117),
				.b5(W2B127),
				.b6(W2B207),
				.b7(W2B217),
				.b8(W2B227),
				.c(c2722B)
);

ninexnine_unit ninexnine_unit_4684(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2B008),
				.b1(W2B018),
				.b2(W2B028),
				.b3(W2B108),
				.b4(W2B118),
				.b5(W2B128),
				.b6(W2B208),
				.b7(W2B218),
				.b8(W2B228),
				.c(c2822B)
);

ninexnine_unit ninexnine_unit_4685(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2B009),
				.b1(W2B019),
				.b2(W2B029),
				.b3(W2B109),
				.b4(W2B119),
				.b5(W2B129),
				.b6(W2B209),
				.b7(W2B219),
				.b8(W2B229),
				.c(c2922B)
);

ninexnine_unit ninexnine_unit_4686(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2B00A),
				.b1(W2B01A),
				.b2(W2B02A),
				.b3(W2B10A),
				.b4(W2B11A),
				.b5(W2B12A),
				.b6(W2B20A),
				.b7(W2B21A),
				.b8(W2B22A),
				.c(c2A22B)
);

ninexnine_unit ninexnine_unit_4687(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2B00B),
				.b1(W2B01B),
				.b2(W2B02B),
				.b3(W2B10B),
				.b4(W2B11B),
				.b5(W2B12B),
				.b6(W2B20B),
				.b7(W2B21B),
				.b8(W2B22B),
				.c(c2B22B)
);

ninexnine_unit ninexnine_unit_4688(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2B00C),
				.b1(W2B01C),
				.b2(W2B02C),
				.b3(W2B10C),
				.b4(W2B11C),
				.b5(W2B12C),
				.b6(W2B20C),
				.b7(W2B21C),
				.b8(W2B22C),
				.c(c2C22B)
);

ninexnine_unit ninexnine_unit_4689(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2B00D),
				.b1(W2B01D),
				.b2(W2B02D),
				.b3(W2B10D),
				.b4(W2B11D),
				.b5(W2B12D),
				.b6(W2B20D),
				.b7(W2B21D),
				.b8(W2B22D),
				.c(c2D22B)
);

ninexnine_unit ninexnine_unit_4690(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2B00E),
				.b1(W2B01E),
				.b2(W2B02E),
				.b3(W2B10E),
				.b4(W2B11E),
				.b5(W2B12E),
				.b6(W2B20E),
				.b7(W2B21E),
				.b8(W2B22E),
				.c(c2E22B)
);

ninexnine_unit ninexnine_unit_4691(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2B00F),
				.b1(W2B01F),
				.b2(W2B02F),
				.b3(W2B10F),
				.b4(W2B11F),
				.b5(W2B12F),
				.b6(W2B20F),
				.b7(W2B21F),
				.b8(W2B22F),
				.c(c2F22B)
);

assign C222B=c2022B+c2122B+c2222B+c2322B+c2422B+c2522B+c2622B+c2722B+c2822B+c2922B+c2A22B+c2B22B+c2C22B+c2D22B+c2E22B+c2F22B;
assign A222B=(C222B>=0)?1:0;

assign P322B=A222B;

ninexnine_unit ninexnine_unit_4692(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2000C)
);

ninexnine_unit ninexnine_unit_4693(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2100C)
);

ninexnine_unit ninexnine_unit_4694(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2200C)
);

ninexnine_unit ninexnine_unit_4695(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2300C)
);

ninexnine_unit ninexnine_unit_4696(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2400C)
);

ninexnine_unit ninexnine_unit_4697(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2500C)
);

ninexnine_unit ninexnine_unit_4698(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2600C)
);

ninexnine_unit ninexnine_unit_4699(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2700C)
);

ninexnine_unit ninexnine_unit_4700(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2C008),
				.b1(W2C018),
				.b2(W2C028),
				.b3(W2C108),
				.b4(W2C118),
				.b5(W2C128),
				.b6(W2C208),
				.b7(W2C218),
				.b8(W2C228),
				.c(c2800C)
);

ninexnine_unit ninexnine_unit_4701(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2C009),
				.b1(W2C019),
				.b2(W2C029),
				.b3(W2C109),
				.b4(W2C119),
				.b5(W2C129),
				.b6(W2C209),
				.b7(W2C219),
				.b8(W2C229),
				.c(c2900C)
);

ninexnine_unit ninexnine_unit_4702(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2C00A),
				.b1(W2C01A),
				.b2(W2C02A),
				.b3(W2C10A),
				.b4(W2C11A),
				.b5(W2C12A),
				.b6(W2C20A),
				.b7(W2C21A),
				.b8(W2C22A),
				.c(c2A00C)
);

ninexnine_unit ninexnine_unit_4703(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2C00B),
				.b1(W2C01B),
				.b2(W2C02B),
				.b3(W2C10B),
				.b4(W2C11B),
				.b5(W2C12B),
				.b6(W2C20B),
				.b7(W2C21B),
				.b8(W2C22B),
				.c(c2B00C)
);

ninexnine_unit ninexnine_unit_4704(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2C00C),
				.b1(W2C01C),
				.b2(W2C02C),
				.b3(W2C10C),
				.b4(W2C11C),
				.b5(W2C12C),
				.b6(W2C20C),
				.b7(W2C21C),
				.b8(W2C22C),
				.c(c2C00C)
);

ninexnine_unit ninexnine_unit_4705(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2C00D),
				.b1(W2C01D),
				.b2(W2C02D),
				.b3(W2C10D),
				.b4(W2C11D),
				.b5(W2C12D),
				.b6(W2C20D),
				.b7(W2C21D),
				.b8(W2C22D),
				.c(c2D00C)
);

ninexnine_unit ninexnine_unit_4706(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2C00E),
				.b1(W2C01E),
				.b2(W2C02E),
				.b3(W2C10E),
				.b4(W2C11E),
				.b5(W2C12E),
				.b6(W2C20E),
				.b7(W2C21E),
				.b8(W2C22E),
				.c(c2E00C)
);

ninexnine_unit ninexnine_unit_4707(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2C00F),
				.b1(W2C01F),
				.b2(W2C02F),
				.b3(W2C10F),
				.b4(W2C11F),
				.b5(W2C12F),
				.b6(W2C20F),
				.b7(W2C21F),
				.b8(W2C22F),
				.c(c2F00C)
);

assign C200C=c2000C+c2100C+c2200C+c2300C+c2400C+c2500C+c2600C+c2700C+c2800C+c2900C+c2A00C+c2B00C+c2C00C+c2D00C+c2E00C+c2F00C;
assign A200C=(C200C>=0)?1:0;

assign P300C=A200C;

ninexnine_unit ninexnine_unit_4708(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2001C)
);

ninexnine_unit ninexnine_unit_4709(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2101C)
);

ninexnine_unit ninexnine_unit_4710(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2201C)
);

ninexnine_unit ninexnine_unit_4711(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2301C)
);

ninexnine_unit ninexnine_unit_4712(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2401C)
);

ninexnine_unit ninexnine_unit_4713(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2501C)
);

ninexnine_unit ninexnine_unit_4714(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2601C)
);

ninexnine_unit ninexnine_unit_4715(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2701C)
);

ninexnine_unit ninexnine_unit_4716(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2C008),
				.b1(W2C018),
				.b2(W2C028),
				.b3(W2C108),
				.b4(W2C118),
				.b5(W2C128),
				.b6(W2C208),
				.b7(W2C218),
				.b8(W2C228),
				.c(c2801C)
);

ninexnine_unit ninexnine_unit_4717(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2C009),
				.b1(W2C019),
				.b2(W2C029),
				.b3(W2C109),
				.b4(W2C119),
				.b5(W2C129),
				.b6(W2C209),
				.b7(W2C219),
				.b8(W2C229),
				.c(c2901C)
);

ninexnine_unit ninexnine_unit_4718(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2C00A),
				.b1(W2C01A),
				.b2(W2C02A),
				.b3(W2C10A),
				.b4(W2C11A),
				.b5(W2C12A),
				.b6(W2C20A),
				.b7(W2C21A),
				.b8(W2C22A),
				.c(c2A01C)
);

ninexnine_unit ninexnine_unit_4719(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2C00B),
				.b1(W2C01B),
				.b2(W2C02B),
				.b3(W2C10B),
				.b4(W2C11B),
				.b5(W2C12B),
				.b6(W2C20B),
				.b7(W2C21B),
				.b8(W2C22B),
				.c(c2B01C)
);

ninexnine_unit ninexnine_unit_4720(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2C00C),
				.b1(W2C01C),
				.b2(W2C02C),
				.b3(W2C10C),
				.b4(W2C11C),
				.b5(W2C12C),
				.b6(W2C20C),
				.b7(W2C21C),
				.b8(W2C22C),
				.c(c2C01C)
);

ninexnine_unit ninexnine_unit_4721(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2C00D),
				.b1(W2C01D),
				.b2(W2C02D),
				.b3(W2C10D),
				.b4(W2C11D),
				.b5(W2C12D),
				.b6(W2C20D),
				.b7(W2C21D),
				.b8(W2C22D),
				.c(c2D01C)
);

ninexnine_unit ninexnine_unit_4722(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2C00E),
				.b1(W2C01E),
				.b2(W2C02E),
				.b3(W2C10E),
				.b4(W2C11E),
				.b5(W2C12E),
				.b6(W2C20E),
				.b7(W2C21E),
				.b8(W2C22E),
				.c(c2E01C)
);

ninexnine_unit ninexnine_unit_4723(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2C00F),
				.b1(W2C01F),
				.b2(W2C02F),
				.b3(W2C10F),
				.b4(W2C11F),
				.b5(W2C12F),
				.b6(W2C20F),
				.b7(W2C21F),
				.b8(W2C22F),
				.c(c2F01C)
);

assign C201C=c2001C+c2101C+c2201C+c2301C+c2401C+c2501C+c2601C+c2701C+c2801C+c2901C+c2A01C+c2B01C+c2C01C+c2D01C+c2E01C+c2F01C;
assign A201C=(C201C>=0)?1:0;

assign P301C=A201C;

ninexnine_unit ninexnine_unit_4724(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2002C)
);

ninexnine_unit ninexnine_unit_4725(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2102C)
);

ninexnine_unit ninexnine_unit_4726(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2202C)
);

ninexnine_unit ninexnine_unit_4727(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2302C)
);

ninexnine_unit ninexnine_unit_4728(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2402C)
);

ninexnine_unit ninexnine_unit_4729(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2502C)
);

ninexnine_unit ninexnine_unit_4730(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2602C)
);

ninexnine_unit ninexnine_unit_4731(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2702C)
);

ninexnine_unit ninexnine_unit_4732(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2C008),
				.b1(W2C018),
				.b2(W2C028),
				.b3(W2C108),
				.b4(W2C118),
				.b5(W2C128),
				.b6(W2C208),
				.b7(W2C218),
				.b8(W2C228),
				.c(c2802C)
);

ninexnine_unit ninexnine_unit_4733(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2C009),
				.b1(W2C019),
				.b2(W2C029),
				.b3(W2C109),
				.b4(W2C119),
				.b5(W2C129),
				.b6(W2C209),
				.b7(W2C219),
				.b8(W2C229),
				.c(c2902C)
);

ninexnine_unit ninexnine_unit_4734(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2C00A),
				.b1(W2C01A),
				.b2(W2C02A),
				.b3(W2C10A),
				.b4(W2C11A),
				.b5(W2C12A),
				.b6(W2C20A),
				.b7(W2C21A),
				.b8(W2C22A),
				.c(c2A02C)
);

ninexnine_unit ninexnine_unit_4735(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2C00B),
				.b1(W2C01B),
				.b2(W2C02B),
				.b3(W2C10B),
				.b4(W2C11B),
				.b5(W2C12B),
				.b6(W2C20B),
				.b7(W2C21B),
				.b8(W2C22B),
				.c(c2B02C)
);

ninexnine_unit ninexnine_unit_4736(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2C00C),
				.b1(W2C01C),
				.b2(W2C02C),
				.b3(W2C10C),
				.b4(W2C11C),
				.b5(W2C12C),
				.b6(W2C20C),
				.b7(W2C21C),
				.b8(W2C22C),
				.c(c2C02C)
);

ninexnine_unit ninexnine_unit_4737(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2C00D),
				.b1(W2C01D),
				.b2(W2C02D),
				.b3(W2C10D),
				.b4(W2C11D),
				.b5(W2C12D),
				.b6(W2C20D),
				.b7(W2C21D),
				.b8(W2C22D),
				.c(c2D02C)
);

ninexnine_unit ninexnine_unit_4738(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2C00E),
				.b1(W2C01E),
				.b2(W2C02E),
				.b3(W2C10E),
				.b4(W2C11E),
				.b5(W2C12E),
				.b6(W2C20E),
				.b7(W2C21E),
				.b8(W2C22E),
				.c(c2E02C)
);

ninexnine_unit ninexnine_unit_4739(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2C00F),
				.b1(W2C01F),
				.b2(W2C02F),
				.b3(W2C10F),
				.b4(W2C11F),
				.b5(W2C12F),
				.b6(W2C20F),
				.b7(W2C21F),
				.b8(W2C22F),
				.c(c2F02C)
);

assign C202C=c2002C+c2102C+c2202C+c2302C+c2402C+c2502C+c2602C+c2702C+c2802C+c2902C+c2A02C+c2B02C+c2C02C+c2D02C+c2E02C+c2F02C;
assign A202C=(C202C>=0)?1:0;

assign P302C=A202C;

ninexnine_unit ninexnine_unit_4740(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2010C)
);

ninexnine_unit ninexnine_unit_4741(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2110C)
);

ninexnine_unit ninexnine_unit_4742(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2210C)
);

ninexnine_unit ninexnine_unit_4743(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2310C)
);

ninexnine_unit ninexnine_unit_4744(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2410C)
);

ninexnine_unit ninexnine_unit_4745(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2510C)
);

ninexnine_unit ninexnine_unit_4746(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2610C)
);

ninexnine_unit ninexnine_unit_4747(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2710C)
);

ninexnine_unit ninexnine_unit_4748(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2C008),
				.b1(W2C018),
				.b2(W2C028),
				.b3(W2C108),
				.b4(W2C118),
				.b5(W2C128),
				.b6(W2C208),
				.b7(W2C218),
				.b8(W2C228),
				.c(c2810C)
);

ninexnine_unit ninexnine_unit_4749(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2C009),
				.b1(W2C019),
				.b2(W2C029),
				.b3(W2C109),
				.b4(W2C119),
				.b5(W2C129),
				.b6(W2C209),
				.b7(W2C219),
				.b8(W2C229),
				.c(c2910C)
);

ninexnine_unit ninexnine_unit_4750(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2C00A),
				.b1(W2C01A),
				.b2(W2C02A),
				.b3(W2C10A),
				.b4(W2C11A),
				.b5(W2C12A),
				.b6(W2C20A),
				.b7(W2C21A),
				.b8(W2C22A),
				.c(c2A10C)
);

ninexnine_unit ninexnine_unit_4751(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2C00B),
				.b1(W2C01B),
				.b2(W2C02B),
				.b3(W2C10B),
				.b4(W2C11B),
				.b5(W2C12B),
				.b6(W2C20B),
				.b7(W2C21B),
				.b8(W2C22B),
				.c(c2B10C)
);

ninexnine_unit ninexnine_unit_4752(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2C00C),
				.b1(W2C01C),
				.b2(W2C02C),
				.b3(W2C10C),
				.b4(W2C11C),
				.b5(W2C12C),
				.b6(W2C20C),
				.b7(W2C21C),
				.b8(W2C22C),
				.c(c2C10C)
);

ninexnine_unit ninexnine_unit_4753(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2C00D),
				.b1(W2C01D),
				.b2(W2C02D),
				.b3(W2C10D),
				.b4(W2C11D),
				.b5(W2C12D),
				.b6(W2C20D),
				.b7(W2C21D),
				.b8(W2C22D),
				.c(c2D10C)
);

ninexnine_unit ninexnine_unit_4754(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2C00E),
				.b1(W2C01E),
				.b2(W2C02E),
				.b3(W2C10E),
				.b4(W2C11E),
				.b5(W2C12E),
				.b6(W2C20E),
				.b7(W2C21E),
				.b8(W2C22E),
				.c(c2E10C)
);

ninexnine_unit ninexnine_unit_4755(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2C00F),
				.b1(W2C01F),
				.b2(W2C02F),
				.b3(W2C10F),
				.b4(W2C11F),
				.b5(W2C12F),
				.b6(W2C20F),
				.b7(W2C21F),
				.b8(W2C22F),
				.c(c2F10C)
);

assign C210C=c2010C+c2110C+c2210C+c2310C+c2410C+c2510C+c2610C+c2710C+c2810C+c2910C+c2A10C+c2B10C+c2C10C+c2D10C+c2E10C+c2F10C;
assign A210C=(C210C>=0)?1:0;

assign P310C=A210C;

ninexnine_unit ninexnine_unit_4756(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2011C)
);

ninexnine_unit ninexnine_unit_4757(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2111C)
);

ninexnine_unit ninexnine_unit_4758(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2211C)
);

ninexnine_unit ninexnine_unit_4759(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2311C)
);

ninexnine_unit ninexnine_unit_4760(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2411C)
);

ninexnine_unit ninexnine_unit_4761(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2511C)
);

ninexnine_unit ninexnine_unit_4762(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2611C)
);

ninexnine_unit ninexnine_unit_4763(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2711C)
);

ninexnine_unit ninexnine_unit_4764(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2C008),
				.b1(W2C018),
				.b2(W2C028),
				.b3(W2C108),
				.b4(W2C118),
				.b5(W2C128),
				.b6(W2C208),
				.b7(W2C218),
				.b8(W2C228),
				.c(c2811C)
);

ninexnine_unit ninexnine_unit_4765(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2C009),
				.b1(W2C019),
				.b2(W2C029),
				.b3(W2C109),
				.b4(W2C119),
				.b5(W2C129),
				.b6(W2C209),
				.b7(W2C219),
				.b8(W2C229),
				.c(c2911C)
);

ninexnine_unit ninexnine_unit_4766(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2C00A),
				.b1(W2C01A),
				.b2(W2C02A),
				.b3(W2C10A),
				.b4(W2C11A),
				.b5(W2C12A),
				.b6(W2C20A),
				.b7(W2C21A),
				.b8(W2C22A),
				.c(c2A11C)
);

ninexnine_unit ninexnine_unit_4767(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2C00B),
				.b1(W2C01B),
				.b2(W2C02B),
				.b3(W2C10B),
				.b4(W2C11B),
				.b5(W2C12B),
				.b6(W2C20B),
				.b7(W2C21B),
				.b8(W2C22B),
				.c(c2B11C)
);

ninexnine_unit ninexnine_unit_4768(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2C00C),
				.b1(W2C01C),
				.b2(W2C02C),
				.b3(W2C10C),
				.b4(W2C11C),
				.b5(W2C12C),
				.b6(W2C20C),
				.b7(W2C21C),
				.b8(W2C22C),
				.c(c2C11C)
);

ninexnine_unit ninexnine_unit_4769(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2C00D),
				.b1(W2C01D),
				.b2(W2C02D),
				.b3(W2C10D),
				.b4(W2C11D),
				.b5(W2C12D),
				.b6(W2C20D),
				.b7(W2C21D),
				.b8(W2C22D),
				.c(c2D11C)
);

ninexnine_unit ninexnine_unit_4770(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2C00E),
				.b1(W2C01E),
				.b2(W2C02E),
				.b3(W2C10E),
				.b4(W2C11E),
				.b5(W2C12E),
				.b6(W2C20E),
				.b7(W2C21E),
				.b8(W2C22E),
				.c(c2E11C)
);

ninexnine_unit ninexnine_unit_4771(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2C00F),
				.b1(W2C01F),
				.b2(W2C02F),
				.b3(W2C10F),
				.b4(W2C11F),
				.b5(W2C12F),
				.b6(W2C20F),
				.b7(W2C21F),
				.b8(W2C22F),
				.c(c2F11C)
);

assign C211C=c2011C+c2111C+c2211C+c2311C+c2411C+c2511C+c2611C+c2711C+c2811C+c2911C+c2A11C+c2B11C+c2C11C+c2D11C+c2E11C+c2F11C;
assign A211C=(C211C>=0)?1:0;

assign P311C=A211C;

ninexnine_unit ninexnine_unit_4772(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2012C)
);

ninexnine_unit ninexnine_unit_4773(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2112C)
);

ninexnine_unit ninexnine_unit_4774(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2212C)
);

ninexnine_unit ninexnine_unit_4775(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2312C)
);

ninexnine_unit ninexnine_unit_4776(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2412C)
);

ninexnine_unit ninexnine_unit_4777(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2512C)
);

ninexnine_unit ninexnine_unit_4778(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2612C)
);

ninexnine_unit ninexnine_unit_4779(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2712C)
);

ninexnine_unit ninexnine_unit_4780(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2C008),
				.b1(W2C018),
				.b2(W2C028),
				.b3(W2C108),
				.b4(W2C118),
				.b5(W2C128),
				.b6(W2C208),
				.b7(W2C218),
				.b8(W2C228),
				.c(c2812C)
);

ninexnine_unit ninexnine_unit_4781(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2C009),
				.b1(W2C019),
				.b2(W2C029),
				.b3(W2C109),
				.b4(W2C119),
				.b5(W2C129),
				.b6(W2C209),
				.b7(W2C219),
				.b8(W2C229),
				.c(c2912C)
);

ninexnine_unit ninexnine_unit_4782(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2C00A),
				.b1(W2C01A),
				.b2(W2C02A),
				.b3(W2C10A),
				.b4(W2C11A),
				.b5(W2C12A),
				.b6(W2C20A),
				.b7(W2C21A),
				.b8(W2C22A),
				.c(c2A12C)
);

ninexnine_unit ninexnine_unit_4783(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2C00B),
				.b1(W2C01B),
				.b2(W2C02B),
				.b3(W2C10B),
				.b4(W2C11B),
				.b5(W2C12B),
				.b6(W2C20B),
				.b7(W2C21B),
				.b8(W2C22B),
				.c(c2B12C)
);

ninexnine_unit ninexnine_unit_4784(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2C00C),
				.b1(W2C01C),
				.b2(W2C02C),
				.b3(W2C10C),
				.b4(W2C11C),
				.b5(W2C12C),
				.b6(W2C20C),
				.b7(W2C21C),
				.b8(W2C22C),
				.c(c2C12C)
);

ninexnine_unit ninexnine_unit_4785(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2C00D),
				.b1(W2C01D),
				.b2(W2C02D),
				.b3(W2C10D),
				.b4(W2C11D),
				.b5(W2C12D),
				.b6(W2C20D),
				.b7(W2C21D),
				.b8(W2C22D),
				.c(c2D12C)
);

ninexnine_unit ninexnine_unit_4786(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2C00E),
				.b1(W2C01E),
				.b2(W2C02E),
				.b3(W2C10E),
				.b4(W2C11E),
				.b5(W2C12E),
				.b6(W2C20E),
				.b7(W2C21E),
				.b8(W2C22E),
				.c(c2E12C)
);

ninexnine_unit ninexnine_unit_4787(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2C00F),
				.b1(W2C01F),
				.b2(W2C02F),
				.b3(W2C10F),
				.b4(W2C11F),
				.b5(W2C12F),
				.b6(W2C20F),
				.b7(W2C21F),
				.b8(W2C22F),
				.c(c2F12C)
);

assign C212C=c2012C+c2112C+c2212C+c2312C+c2412C+c2512C+c2612C+c2712C+c2812C+c2912C+c2A12C+c2B12C+c2C12C+c2D12C+c2E12C+c2F12C;
assign A212C=(C212C>=0)?1:0;

assign P312C=A212C;

ninexnine_unit ninexnine_unit_4788(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2020C)
);

ninexnine_unit ninexnine_unit_4789(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2120C)
);

ninexnine_unit ninexnine_unit_4790(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2220C)
);

ninexnine_unit ninexnine_unit_4791(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2320C)
);

ninexnine_unit ninexnine_unit_4792(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2420C)
);

ninexnine_unit ninexnine_unit_4793(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2520C)
);

ninexnine_unit ninexnine_unit_4794(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2620C)
);

ninexnine_unit ninexnine_unit_4795(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2720C)
);

ninexnine_unit ninexnine_unit_4796(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2C008),
				.b1(W2C018),
				.b2(W2C028),
				.b3(W2C108),
				.b4(W2C118),
				.b5(W2C128),
				.b6(W2C208),
				.b7(W2C218),
				.b8(W2C228),
				.c(c2820C)
);

ninexnine_unit ninexnine_unit_4797(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2C009),
				.b1(W2C019),
				.b2(W2C029),
				.b3(W2C109),
				.b4(W2C119),
				.b5(W2C129),
				.b6(W2C209),
				.b7(W2C219),
				.b8(W2C229),
				.c(c2920C)
);

ninexnine_unit ninexnine_unit_4798(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2C00A),
				.b1(W2C01A),
				.b2(W2C02A),
				.b3(W2C10A),
				.b4(W2C11A),
				.b5(W2C12A),
				.b6(W2C20A),
				.b7(W2C21A),
				.b8(W2C22A),
				.c(c2A20C)
);

ninexnine_unit ninexnine_unit_4799(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2C00B),
				.b1(W2C01B),
				.b2(W2C02B),
				.b3(W2C10B),
				.b4(W2C11B),
				.b5(W2C12B),
				.b6(W2C20B),
				.b7(W2C21B),
				.b8(W2C22B),
				.c(c2B20C)
);

ninexnine_unit ninexnine_unit_4800(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2C00C),
				.b1(W2C01C),
				.b2(W2C02C),
				.b3(W2C10C),
				.b4(W2C11C),
				.b5(W2C12C),
				.b6(W2C20C),
				.b7(W2C21C),
				.b8(W2C22C),
				.c(c2C20C)
);

ninexnine_unit ninexnine_unit_4801(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2C00D),
				.b1(W2C01D),
				.b2(W2C02D),
				.b3(W2C10D),
				.b4(W2C11D),
				.b5(W2C12D),
				.b6(W2C20D),
				.b7(W2C21D),
				.b8(W2C22D),
				.c(c2D20C)
);

ninexnine_unit ninexnine_unit_4802(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2C00E),
				.b1(W2C01E),
				.b2(W2C02E),
				.b3(W2C10E),
				.b4(W2C11E),
				.b5(W2C12E),
				.b6(W2C20E),
				.b7(W2C21E),
				.b8(W2C22E),
				.c(c2E20C)
);

ninexnine_unit ninexnine_unit_4803(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2C00F),
				.b1(W2C01F),
				.b2(W2C02F),
				.b3(W2C10F),
				.b4(W2C11F),
				.b5(W2C12F),
				.b6(W2C20F),
				.b7(W2C21F),
				.b8(W2C22F),
				.c(c2F20C)
);

assign C220C=c2020C+c2120C+c2220C+c2320C+c2420C+c2520C+c2620C+c2720C+c2820C+c2920C+c2A20C+c2B20C+c2C20C+c2D20C+c2E20C+c2F20C;
assign A220C=(C220C>=0)?1:0;

assign P320C=A220C;

ninexnine_unit ninexnine_unit_4804(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2021C)
);

ninexnine_unit ninexnine_unit_4805(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2121C)
);

ninexnine_unit ninexnine_unit_4806(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2221C)
);

ninexnine_unit ninexnine_unit_4807(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2321C)
);

ninexnine_unit ninexnine_unit_4808(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2421C)
);

ninexnine_unit ninexnine_unit_4809(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2521C)
);

ninexnine_unit ninexnine_unit_4810(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2621C)
);

ninexnine_unit ninexnine_unit_4811(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2721C)
);

ninexnine_unit ninexnine_unit_4812(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2C008),
				.b1(W2C018),
				.b2(W2C028),
				.b3(W2C108),
				.b4(W2C118),
				.b5(W2C128),
				.b6(W2C208),
				.b7(W2C218),
				.b8(W2C228),
				.c(c2821C)
);

ninexnine_unit ninexnine_unit_4813(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2C009),
				.b1(W2C019),
				.b2(W2C029),
				.b3(W2C109),
				.b4(W2C119),
				.b5(W2C129),
				.b6(W2C209),
				.b7(W2C219),
				.b8(W2C229),
				.c(c2921C)
);

ninexnine_unit ninexnine_unit_4814(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2C00A),
				.b1(W2C01A),
				.b2(W2C02A),
				.b3(W2C10A),
				.b4(W2C11A),
				.b5(W2C12A),
				.b6(W2C20A),
				.b7(W2C21A),
				.b8(W2C22A),
				.c(c2A21C)
);

ninexnine_unit ninexnine_unit_4815(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2C00B),
				.b1(W2C01B),
				.b2(W2C02B),
				.b3(W2C10B),
				.b4(W2C11B),
				.b5(W2C12B),
				.b6(W2C20B),
				.b7(W2C21B),
				.b8(W2C22B),
				.c(c2B21C)
);

ninexnine_unit ninexnine_unit_4816(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2C00C),
				.b1(W2C01C),
				.b2(W2C02C),
				.b3(W2C10C),
				.b4(W2C11C),
				.b5(W2C12C),
				.b6(W2C20C),
				.b7(W2C21C),
				.b8(W2C22C),
				.c(c2C21C)
);

ninexnine_unit ninexnine_unit_4817(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2C00D),
				.b1(W2C01D),
				.b2(W2C02D),
				.b3(W2C10D),
				.b4(W2C11D),
				.b5(W2C12D),
				.b6(W2C20D),
				.b7(W2C21D),
				.b8(W2C22D),
				.c(c2D21C)
);

ninexnine_unit ninexnine_unit_4818(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2C00E),
				.b1(W2C01E),
				.b2(W2C02E),
				.b3(W2C10E),
				.b4(W2C11E),
				.b5(W2C12E),
				.b6(W2C20E),
				.b7(W2C21E),
				.b8(W2C22E),
				.c(c2E21C)
);

ninexnine_unit ninexnine_unit_4819(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2C00F),
				.b1(W2C01F),
				.b2(W2C02F),
				.b3(W2C10F),
				.b4(W2C11F),
				.b5(W2C12F),
				.b6(W2C20F),
				.b7(W2C21F),
				.b8(W2C22F),
				.c(c2F21C)
);

assign C221C=c2021C+c2121C+c2221C+c2321C+c2421C+c2521C+c2621C+c2721C+c2821C+c2921C+c2A21C+c2B21C+c2C21C+c2D21C+c2E21C+c2F21C;
assign A221C=(C221C>=0)?1:0;

assign P321C=A221C;

ninexnine_unit ninexnine_unit_4820(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2C000),
				.b1(W2C010),
				.b2(W2C020),
				.b3(W2C100),
				.b4(W2C110),
				.b5(W2C120),
				.b6(W2C200),
				.b7(W2C210),
				.b8(W2C220),
				.c(c2022C)
);

ninexnine_unit ninexnine_unit_4821(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2C001),
				.b1(W2C011),
				.b2(W2C021),
				.b3(W2C101),
				.b4(W2C111),
				.b5(W2C121),
				.b6(W2C201),
				.b7(W2C211),
				.b8(W2C221),
				.c(c2122C)
);

ninexnine_unit ninexnine_unit_4822(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2C002),
				.b1(W2C012),
				.b2(W2C022),
				.b3(W2C102),
				.b4(W2C112),
				.b5(W2C122),
				.b6(W2C202),
				.b7(W2C212),
				.b8(W2C222),
				.c(c2222C)
);

ninexnine_unit ninexnine_unit_4823(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2C003),
				.b1(W2C013),
				.b2(W2C023),
				.b3(W2C103),
				.b4(W2C113),
				.b5(W2C123),
				.b6(W2C203),
				.b7(W2C213),
				.b8(W2C223),
				.c(c2322C)
);

ninexnine_unit ninexnine_unit_4824(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2C004),
				.b1(W2C014),
				.b2(W2C024),
				.b3(W2C104),
				.b4(W2C114),
				.b5(W2C124),
				.b6(W2C204),
				.b7(W2C214),
				.b8(W2C224),
				.c(c2422C)
);

ninexnine_unit ninexnine_unit_4825(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2C005),
				.b1(W2C015),
				.b2(W2C025),
				.b3(W2C105),
				.b4(W2C115),
				.b5(W2C125),
				.b6(W2C205),
				.b7(W2C215),
				.b8(W2C225),
				.c(c2522C)
);

ninexnine_unit ninexnine_unit_4826(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2C006),
				.b1(W2C016),
				.b2(W2C026),
				.b3(W2C106),
				.b4(W2C116),
				.b5(W2C126),
				.b6(W2C206),
				.b7(W2C216),
				.b8(W2C226),
				.c(c2622C)
);

ninexnine_unit ninexnine_unit_4827(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2C007),
				.b1(W2C017),
				.b2(W2C027),
				.b3(W2C107),
				.b4(W2C117),
				.b5(W2C127),
				.b6(W2C207),
				.b7(W2C217),
				.b8(W2C227),
				.c(c2722C)
);

ninexnine_unit ninexnine_unit_4828(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2C008),
				.b1(W2C018),
				.b2(W2C028),
				.b3(W2C108),
				.b4(W2C118),
				.b5(W2C128),
				.b6(W2C208),
				.b7(W2C218),
				.b8(W2C228),
				.c(c2822C)
);

ninexnine_unit ninexnine_unit_4829(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2C009),
				.b1(W2C019),
				.b2(W2C029),
				.b3(W2C109),
				.b4(W2C119),
				.b5(W2C129),
				.b6(W2C209),
				.b7(W2C219),
				.b8(W2C229),
				.c(c2922C)
);

ninexnine_unit ninexnine_unit_4830(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2C00A),
				.b1(W2C01A),
				.b2(W2C02A),
				.b3(W2C10A),
				.b4(W2C11A),
				.b5(W2C12A),
				.b6(W2C20A),
				.b7(W2C21A),
				.b8(W2C22A),
				.c(c2A22C)
);

ninexnine_unit ninexnine_unit_4831(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2C00B),
				.b1(W2C01B),
				.b2(W2C02B),
				.b3(W2C10B),
				.b4(W2C11B),
				.b5(W2C12B),
				.b6(W2C20B),
				.b7(W2C21B),
				.b8(W2C22B),
				.c(c2B22C)
);

ninexnine_unit ninexnine_unit_4832(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2C00C),
				.b1(W2C01C),
				.b2(W2C02C),
				.b3(W2C10C),
				.b4(W2C11C),
				.b5(W2C12C),
				.b6(W2C20C),
				.b7(W2C21C),
				.b8(W2C22C),
				.c(c2C22C)
);

ninexnine_unit ninexnine_unit_4833(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2C00D),
				.b1(W2C01D),
				.b2(W2C02D),
				.b3(W2C10D),
				.b4(W2C11D),
				.b5(W2C12D),
				.b6(W2C20D),
				.b7(W2C21D),
				.b8(W2C22D),
				.c(c2D22C)
);

ninexnine_unit ninexnine_unit_4834(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2C00E),
				.b1(W2C01E),
				.b2(W2C02E),
				.b3(W2C10E),
				.b4(W2C11E),
				.b5(W2C12E),
				.b6(W2C20E),
				.b7(W2C21E),
				.b8(W2C22E),
				.c(c2E22C)
);

ninexnine_unit ninexnine_unit_4835(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2C00F),
				.b1(W2C01F),
				.b2(W2C02F),
				.b3(W2C10F),
				.b4(W2C11F),
				.b5(W2C12F),
				.b6(W2C20F),
				.b7(W2C21F),
				.b8(W2C22F),
				.c(c2F22C)
);

assign C222C=c2022C+c2122C+c2222C+c2322C+c2422C+c2522C+c2622C+c2722C+c2822C+c2922C+c2A22C+c2B22C+c2C22C+c2D22C+c2E22C+c2F22C;
assign A222C=(C222C>=0)?1:0;

assign P322C=A222C;

ninexnine_unit ninexnine_unit_4836(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2000D)
);

ninexnine_unit ninexnine_unit_4837(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2100D)
);

ninexnine_unit ninexnine_unit_4838(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2200D)
);

ninexnine_unit ninexnine_unit_4839(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2300D)
);

ninexnine_unit ninexnine_unit_4840(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2400D)
);

ninexnine_unit ninexnine_unit_4841(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2500D)
);

ninexnine_unit ninexnine_unit_4842(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2600D)
);

ninexnine_unit ninexnine_unit_4843(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2700D)
);

ninexnine_unit ninexnine_unit_4844(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2D008),
				.b1(W2D018),
				.b2(W2D028),
				.b3(W2D108),
				.b4(W2D118),
				.b5(W2D128),
				.b6(W2D208),
				.b7(W2D218),
				.b8(W2D228),
				.c(c2800D)
);

ninexnine_unit ninexnine_unit_4845(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2D009),
				.b1(W2D019),
				.b2(W2D029),
				.b3(W2D109),
				.b4(W2D119),
				.b5(W2D129),
				.b6(W2D209),
				.b7(W2D219),
				.b8(W2D229),
				.c(c2900D)
);

ninexnine_unit ninexnine_unit_4846(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2D00A),
				.b1(W2D01A),
				.b2(W2D02A),
				.b3(W2D10A),
				.b4(W2D11A),
				.b5(W2D12A),
				.b6(W2D20A),
				.b7(W2D21A),
				.b8(W2D22A),
				.c(c2A00D)
);

ninexnine_unit ninexnine_unit_4847(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2D00B),
				.b1(W2D01B),
				.b2(W2D02B),
				.b3(W2D10B),
				.b4(W2D11B),
				.b5(W2D12B),
				.b6(W2D20B),
				.b7(W2D21B),
				.b8(W2D22B),
				.c(c2B00D)
);

ninexnine_unit ninexnine_unit_4848(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2D00C),
				.b1(W2D01C),
				.b2(W2D02C),
				.b3(W2D10C),
				.b4(W2D11C),
				.b5(W2D12C),
				.b6(W2D20C),
				.b7(W2D21C),
				.b8(W2D22C),
				.c(c2C00D)
);

ninexnine_unit ninexnine_unit_4849(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2D00D),
				.b1(W2D01D),
				.b2(W2D02D),
				.b3(W2D10D),
				.b4(W2D11D),
				.b5(W2D12D),
				.b6(W2D20D),
				.b7(W2D21D),
				.b8(W2D22D),
				.c(c2D00D)
);

ninexnine_unit ninexnine_unit_4850(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2D00E),
				.b1(W2D01E),
				.b2(W2D02E),
				.b3(W2D10E),
				.b4(W2D11E),
				.b5(W2D12E),
				.b6(W2D20E),
				.b7(W2D21E),
				.b8(W2D22E),
				.c(c2E00D)
);

ninexnine_unit ninexnine_unit_4851(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2D00F),
				.b1(W2D01F),
				.b2(W2D02F),
				.b3(W2D10F),
				.b4(W2D11F),
				.b5(W2D12F),
				.b6(W2D20F),
				.b7(W2D21F),
				.b8(W2D22F),
				.c(c2F00D)
);

assign C200D=c2000D+c2100D+c2200D+c2300D+c2400D+c2500D+c2600D+c2700D+c2800D+c2900D+c2A00D+c2B00D+c2C00D+c2D00D+c2E00D+c2F00D;
assign A200D=(C200D>=0)?1:0;

assign P300D=A200D;

ninexnine_unit ninexnine_unit_4852(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2001D)
);

ninexnine_unit ninexnine_unit_4853(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2101D)
);

ninexnine_unit ninexnine_unit_4854(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2201D)
);

ninexnine_unit ninexnine_unit_4855(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2301D)
);

ninexnine_unit ninexnine_unit_4856(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2401D)
);

ninexnine_unit ninexnine_unit_4857(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2501D)
);

ninexnine_unit ninexnine_unit_4858(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2601D)
);

ninexnine_unit ninexnine_unit_4859(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2701D)
);

ninexnine_unit ninexnine_unit_4860(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2D008),
				.b1(W2D018),
				.b2(W2D028),
				.b3(W2D108),
				.b4(W2D118),
				.b5(W2D128),
				.b6(W2D208),
				.b7(W2D218),
				.b8(W2D228),
				.c(c2801D)
);

ninexnine_unit ninexnine_unit_4861(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2D009),
				.b1(W2D019),
				.b2(W2D029),
				.b3(W2D109),
				.b4(W2D119),
				.b5(W2D129),
				.b6(W2D209),
				.b7(W2D219),
				.b8(W2D229),
				.c(c2901D)
);

ninexnine_unit ninexnine_unit_4862(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2D00A),
				.b1(W2D01A),
				.b2(W2D02A),
				.b3(W2D10A),
				.b4(W2D11A),
				.b5(W2D12A),
				.b6(W2D20A),
				.b7(W2D21A),
				.b8(W2D22A),
				.c(c2A01D)
);

ninexnine_unit ninexnine_unit_4863(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2D00B),
				.b1(W2D01B),
				.b2(W2D02B),
				.b3(W2D10B),
				.b4(W2D11B),
				.b5(W2D12B),
				.b6(W2D20B),
				.b7(W2D21B),
				.b8(W2D22B),
				.c(c2B01D)
);

ninexnine_unit ninexnine_unit_4864(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2D00C),
				.b1(W2D01C),
				.b2(W2D02C),
				.b3(W2D10C),
				.b4(W2D11C),
				.b5(W2D12C),
				.b6(W2D20C),
				.b7(W2D21C),
				.b8(W2D22C),
				.c(c2C01D)
);

ninexnine_unit ninexnine_unit_4865(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2D00D),
				.b1(W2D01D),
				.b2(W2D02D),
				.b3(W2D10D),
				.b4(W2D11D),
				.b5(W2D12D),
				.b6(W2D20D),
				.b7(W2D21D),
				.b8(W2D22D),
				.c(c2D01D)
);

ninexnine_unit ninexnine_unit_4866(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2D00E),
				.b1(W2D01E),
				.b2(W2D02E),
				.b3(W2D10E),
				.b4(W2D11E),
				.b5(W2D12E),
				.b6(W2D20E),
				.b7(W2D21E),
				.b8(W2D22E),
				.c(c2E01D)
);

ninexnine_unit ninexnine_unit_4867(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2D00F),
				.b1(W2D01F),
				.b2(W2D02F),
				.b3(W2D10F),
				.b4(W2D11F),
				.b5(W2D12F),
				.b6(W2D20F),
				.b7(W2D21F),
				.b8(W2D22F),
				.c(c2F01D)
);

assign C201D=c2001D+c2101D+c2201D+c2301D+c2401D+c2501D+c2601D+c2701D+c2801D+c2901D+c2A01D+c2B01D+c2C01D+c2D01D+c2E01D+c2F01D;
assign A201D=(C201D>=0)?1:0;

assign P301D=A201D;

ninexnine_unit ninexnine_unit_4868(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2002D)
);

ninexnine_unit ninexnine_unit_4869(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2102D)
);

ninexnine_unit ninexnine_unit_4870(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2202D)
);

ninexnine_unit ninexnine_unit_4871(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2302D)
);

ninexnine_unit ninexnine_unit_4872(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2402D)
);

ninexnine_unit ninexnine_unit_4873(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2502D)
);

ninexnine_unit ninexnine_unit_4874(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2602D)
);

ninexnine_unit ninexnine_unit_4875(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2702D)
);

ninexnine_unit ninexnine_unit_4876(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2D008),
				.b1(W2D018),
				.b2(W2D028),
				.b3(W2D108),
				.b4(W2D118),
				.b5(W2D128),
				.b6(W2D208),
				.b7(W2D218),
				.b8(W2D228),
				.c(c2802D)
);

ninexnine_unit ninexnine_unit_4877(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2D009),
				.b1(W2D019),
				.b2(W2D029),
				.b3(W2D109),
				.b4(W2D119),
				.b5(W2D129),
				.b6(W2D209),
				.b7(W2D219),
				.b8(W2D229),
				.c(c2902D)
);

ninexnine_unit ninexnine_unit_4878(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2D00A),
				.b1(W2D01A),
				.b2(W2D02A),
				.b3(W2D10A),
				.b4(W2D11A),
				.b5(W2D12A),
				.b6(W2D20A),
				.b7(W2D21A),
				.b8(W2D22A),
				.c(c2A02D)
);

ninexnine_unit ninexnine_unit_4879(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2D00B),
				.b1(W2D01B),
				.b2(W2D02B),
				.b3(W2D10B),
				.b4(W2D11B),
				.b5(W2D12B),
				.b6(W2D20B),
				.b7(W2D21B),
				.b8(W2D22B),
				.c(c2B02D)
);

ninexnine_unit ninexnine_unit_4880(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2D00C),
				.b1(W2D01C),
				.b2(W2D02C),
				.b3(W2D10C),
				.b4(W2D11C),
				.b5(W2D12C),
				.b6(W2D20C),
				.b7(W2D21C),
				.b8(W2D22C),
				.c(c2C02D)
);

ninexnine_unit ninexnine_unit_4881(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2D00D),
				.b1(W2D01D),
				.b2(W2D02D),
				.b3(W2D10D),
				.b4(W2D11D),
				.b5(W2D12D),
				.b6(W2D20D),
				.b7(W2D21D),
				.b8(W2D22D),
				.c(c2D02D)
);

ninexnine_unit ninexnine_unit_4882(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2D00E),
				.b1(W2D01E),
				.b2(W2D02E),
				.b3(W2D10E),
				.b4(W2D11E),
				.b5(W2D12E),
				.b6(W2D20E),
				.b7(W2D21E),
				.b8(W2D22E),
				.c(c2E02D)
);

ninexnine_unit ninexnine_unit_4883(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2D00F),
				.b1(W2D01F),
				.b2(W2D02F),
				.b3(W2D10F),
				.b4(W2D11F),
				.b5(W2D12F),
				.b6(W2D20F),
				.b7(W2D21F),
				.b8(W2D22F),
				.c(c2F02D)
);

assign C202D=c2002D+c2102D+c2202D+c2302D+c2402D+c2502D+c2602D+c2702D+c2802D+c2902D+c2A02D+c2B02D+c2C02D+c2D02D+c2E02D+c2F02D;
assign A202D=(C202D>=0)?1:0;

assign P302D=A202D;

ninexnine_unit ninexnine_unit_4884(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2010D)
);

ninexnine_unit ninexnine_unit_4885(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2110D)
);

ninexnine_unit ninexnine_unit_4886(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2210D)
);

ninexnine_unit ninexnine_unit_4887(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2310D)
);

ninexnine_unit ninexnine_unit_4888(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2410D)
);

ninexnine_unit ninexnine_unit_4889(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2510D)
);

ninexnine_unit ninexnine_unit_4890(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2610D)
);

ninexnine_unit ninexnine_unit_4891(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2710D)
);

ninexnine_unit ninexnine_unit_4892(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2D008),
				.b1(W2D018),
				.b2(W2D028),
				.b3(W2D108),
				.b4(W2D118),
				.b5(W2D128),
				.b6(W2D208),
				.b7(W2D218),
				.b8(W2D228),
				.c(c2810D)
);

ninexnine_unit ninexnine_unit_4893(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2D009),
				.b1(W2D019),
				.b2(W2D029),
				.b3(W2D109),
				.b4(W2D119),
				.b5(W2D129),
				.b6(W2D209),
				.b7(W2D219),
				.b8(W2D229),
				.c(c2910D)
);

ninexnine_unit ninexnine_unit_4894(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2D00A),
				.b1(W2D01A),
				.b2(W2D02A),
				.b3(W2D10A),
				.b4(W2D11A),
				.b5(W2D12A),
				.b6(W2D20A),
				.b7(W2D21A),
				.b8(W2D22A),
				.c(c2A10D)
);

ninexnine_unit ninexnine_unit_4895(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2D00B),
				.b1(W2D01B),
				.b2(W2D02B),
				.b3(W2D10B),
				.b4(W2D11B),
				.b5(W2D12B),
				.b6(W2D20B),
				.b7(W2D21B),
				.b8(W2D22B),
				.c(c2B10D)
);

ninexnine_unit ninexnine_unit_4896(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2D00C),
				.b1(W2D01C),
				.b2(W2D02C),
				.b3(W2D10C),
				.b4(W2D11C),
				.b5(W2D12C),
				.b6(W2D20C),
				.b7(W2D21C),
				.b8(W2D22C),
				.c(c2C10D)
);

ninexnine_unit ninexnine_unit_4897(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2D00D),
				.b1(W2D01D),
				.b2(W2D02D),
				.b3(W2D10D),
				.b4(W2D11D),
				.b5(W2D12D),
				.b6(W2D20D),
				.b7(W2D21D),
				.b8(W2D22D),
				.c(c2D10D)
);

ninexnine_unit ninexnine_unit_4898(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2D00E),
				.b1(W2D01E),
				.b2(W2D02E),
				.b3(W2D10E),
				.b4(W2D11E),
				.b5(W2D12E),
				.b6(W2D20E),
				.b7(W2D21E),
				.b8(W2D22E),
				.c(c2E10D)
);

ninexnine_unit ninexnine_unit_4899(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2D00F),
				.b1(W2D01F),
				.b2(W2D02F),
				.b3(W2D10F),
				.b4(W2D11F),
				.b5(W2D12F),
				.b6(W2D20F),
				.b7(W2D21F),
				.b8(W2D22F),
				.c(c2F10D)
);

assign C210D=c2010D+c2110D+c2210D+c2310D+c2410D+c2510D+c2610D+c2710D+c2810D+c2910D+c2A10D+c2B10D+c2C10D+c2D10D+c2E10D+c2F10D;
assign A210D=(C210D>=0)?1:0;

assign P310D=A210D;

ninexnine_unit ninexnine_unit_4900(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2011D)
);

ninexnine_unit ninexnine_unit_4901(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2111D)
);

ninexnine_unit ninexnine_unit_4902(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2211D)
);

ninexnine_unit ninexnine_unit_4903(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2311D)
);

ninexnine_unit ninexnine_unit_4904(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2411D)
);

ninexnine_unit ninexnine_unit_4905(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2511D)
);

ninexnine_unit ninexnine_unit_4906(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2611D)
);

ninexnine_unit ninexnine_unit_4907(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2711D)
);

ninexnine_unit ninexnine_unit_4908(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2D008),
				.b1(W2D018),
				.b2(W2D028),
				.b3(W2D108),
				.b4(W2D118),
				.b5(W2D128),
				.b6(W2D208),
				.b7(W2D218),
				.b8(W2D228),
				.c(c2811D)
);

ninexnine_unit ninexnine_unit_4909(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2D009),
				.b1(W2D019),
				.b2(W2D029),
				.b3(W2D109),
				.b4(W2D119),
				.b5(W2D129),
				.b6(W2D209),
				.b7(W2D219),
				.b8(W2D229),
				.c(c2911D)
);

ninexnine_unit ninexnine_unit_4910(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2D00A),
				.b1(W2D01A),
				.b2(W2D02A),
				.b3(W2D10A),
				.b4(W2D11A),
				.b5(W2D12A),
				.b6(W2D20A),
				.b7(W2D21A),
				.b8(W2D22A),
				.c(c2A11D)
);

ninexnine_unit ninexnine_unit_4911(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2D00B),
				.b1(W2D01B),
				.b2(W2D02B),
				.b3(W2D10B),
				.b4(W2D11B),
				.b5(W2D12B),
				.b6(W2D20B),
				.b7(W2D21B),
				.b8(W2D22B),
				.c(c2B11D)
);

ninexnine_unit ninexnine_unit_4912(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2D00C),
				.b1(W2D01C),
				.b2(W2D02C),
				.b3(W2D10C),
				.b4(W2D11C),
				.b5(W2D12C),
				.b6(W2D20C),
				.b7(W2D21C),
				.b8(W2D22C),
				.c(c2C11D)
);

ninexnine_unit ninexnine_unit_4913(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2D00D),
				.b1(W2D01D),
				.b2(W2D02D),
				.b3(W2D10D),
				.b4(W2D11D),
				.b5(W2D12D),
				.b6(W2D20D),
				.b7(W2D21D),
				.b8(W2D22D),
				.c(c2D11D)
);

ninexnine_unit ninexnine_unit_4914(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2D00E),
				.b1(W2D01E),
				.b2(W2D02E),
				.b3(W2D10E),
				.b4(W2D11E),
				.b5(W2D12E),
				.b6(W2D20E),
				.b7(W2D21E),
				.b8(W2D22E),
				.c(c2E11D)
);

ninexnine_unit ninexnine_unit_4915(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2D00F),
				.b1(W2D01F),
				.b2(W2D02F),
				.b3(W2D10F),
				.b4(W2D11F),
				.b5(W2D12F),
				.b6(W2D20F),
				.b7(W2D21F),
				.b8(W2D22F),
				.c(c2F11D)
);

assign C211D=c2011D+c2111D+c2211D+c2311D+c2411D+c2511D+c2611D+c2711D+c2811D+c2911D+c2A11D+c2B11D+c2C11D+c2D11D+c2E11D+c2F11D;
assign A211D=(C211D>=0)?1:0;

assign P311D=A211D;

ninexnine_unit ninexnine_unit_4916(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2012D)
);

ninexnine_unit ninexnine_unit_4917(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2112D)
);

ninexnine_unit ninexnine_unit_4918(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2212D)
);

ninexnine_unit ninexnine_unit_4919(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2312D)
);

ninexnine_unit ninexnine_unit_4920(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2412D)
);

ninexnine_unit ninexnine_unit_4921(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2512D)
);

ninexnine_unit ninexnine_unit_4922(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2612D)
);

ninexnine_unit ninexnine_unit_4923(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2712D)
);

ninexnine_unit ninexnine_unit_4924(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2D008),
				.b1(W2D018),
				.b2(W2D028),
				.b3(W2D108),
				.b4(W2D118),
				.b5(W2D128),
				.b6(W2D208),
				.b7(W2D218),
				.b8(W2D228),
				.c(c2812D)
);

ninexnine_unit ninexnine_unit_4925(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2D009),
				.b1(W2D019),
				.b2(W2D029),
				.b3(W2D109),
				.b4(W2D119),
				.b5(W2D129),
				.b6(W2D209),
				.b7(W2D219),
				.b8(W2D229),
				.c(c2912D)
);

ninexnine_unit ninexnine_unit_4926(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2D00A),
				.b1(W2D01A),
				.b2(W2D02A),
				.b3(W2D10A),
				.b4(W2D11A),
				.b5(W2D12A),
				.b6(W2D20A),
				.b7(W2D21A),
				.b8(W2D22A),
				.c(c2A12D)
);

ninexnine_unit ninexnine_unit_4927(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2D00B),
				.b1(W2D01B),
				.b2(W2D02B),
				.b3(W2D10B),
				.b4(W2D11B),
				.b5(W2D12B),
				.b6(W2D20B),
				.b7(W2D21B),
				.b8(W2D22B),
				.c(c2B12D)
);

ninexnine_unit ninexnine_unit_4928(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2D00C),
				.b1(W2D01C),
				.b2(W2D02C),
				.b3(W2D10C),
				.b4(W2D11C),
				.b5(W2D12C),
				.b6(W2D20C),
				.b7(W2D21C),
				.b8(W2D22C),
				.c(c2C12D)
);

ninexnine_unit ninexnine_unit_4929(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2D00D),
				.b1(W2D01D),
				.b2(W2D02D),
				.b3(W2D10D),
				.b4(W2D11D),
				.b5(W2D12D),
				.b6(W2D20D),
				.b7(W2D21D),
				.b8(W2D22D),
				.c(c2D12D)
);

ninexnine_unit ninexnine_unit_4930(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2D00E),
				.b1(W2D01E),
				.b2(W2D02E),
				.b3(W2D10E),
				.b4(W2D11E),
				.b5(W2D12E),
				.b6(W2D20E),
				.b7(W2D21E),
				.b8(W2D22E),
				.c(c2E12D)
);

ninexnine_unit ninexnine_unit_4931(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2D00F),
				.b1(W2D01F),
				.b2(W2D02F),
				.b3(W2D10F),
				.b4(W2D11F),
				.b5(W2D12F),
				.b6(W2D20F),
				.b7(W2D21F),
				.b8(W2D22F),
				.c(c2F12D)
);

assign C212D=c2012D+c2112D+c2212D+c2312D+c2412D+c2512D+c2612D+c2712D+c2812D+c2912D+c2A12D+c2B12D+c2C12D+c2D12D+c2E12D+c2F12D;
assign A212D=(C212D>=0)?1:0;

assign P312D=A212D;

ninexnine_unit ninexnine_unit_4932(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2020D)
);

ninexnine_unit ninexnine_unit_4933(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2120D)
);

ninexnine_unit ninexnine_unit_4934(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2220D)
);

ninexnine_unit ninexnine_unit_4935(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2320D)
);

ninexnine_unit ninexnine_unit_4936(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2420D)
);

ninexnine_unit ninexnine_unit_4937(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2520D)
);

ninexnine_unit ninexnine_unit_4938(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2620D)
);

ninexnine_unit ninexnine_unit_4939(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2720D)
);

ninexnine_unit ninexnine_unit_4940(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2D008),
				.b1(W2D018),
				.b2(W2D028),
				.b3(W2D108),
				.b4(W2D118),
				.b5(W2D128),
				.b6(W2D208),
				.b7(W2D218),
				.b8(W2D228),
				.c(c2820D)
);

ninexnine_unit ninexnine_unit_4941(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2D009),
				.b1(W2D019),
				.b2(W2D029),
				.b3(W2D109),
				.b4(W2D119),
				.b5(W2D129),
				.b6(W2D209),
				.b7(W2D219),
				.b8(W2D229),
				.c(c2920D)
);

ninexnine_unit ninexnine_unit_4942(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2D00A),
				.b1(W2D01A),
				.b2(W2D02A),
				.b3(W2D10A),
				.b4(W2D11A),
				.b5(W2D12A),
				.b6(W2D20A),
				.b7(W2D21A),
				.b8(W2D22A),
				.c(c2A20D)
);

ninexnine_unit ninexnine_unit_4943(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2D00B),
				.b1(W2D01B),
				.b2(W2D02B),
				.b3(W2D10B),
				.b4(W2D11B),
				.b5(W2D12B),
				.b6(W2D20B),
				.b7(W2D21B),
				.b8(W2D22B),
				.c(c2B20D)
);

ninexnine_unit ninexnine_unit_4944(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2D00C),
				.b1(W2D01C),
				.b2(W2D02C),
				.b3(W2D10C),
				.b4(W2D11C),
				.b5(W2D12C),
				.b6(W2D20C),
				.b7(W2D21C),
				.b8(W2D22C),
				.c(c2C20D)
);

ninexnine_unit ninexnine_unit_4945(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2D00D),
				.b1(W2D01D),
				.b2(W2D02D),
				.b3(W2D10D),
				.b4(W2D11D),
				.b5(W2D12D),
				.b6(W2D20D),
				.b7(W2D21D),
				.b8(W2D22D),
				.c(c2D20D)
);

ninexnine_unit ninexnine_unit_4946(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2D00E),
				.b1(W2D01E),
				.b2(W2D02E),
				.b3(W2D10E),
				.b4(W2D11E),
				.b5(W2D12E),
				.b6(W2D20E),
				.b7(W2D21E),
				.b8(W2D22E),
				.c(c2E20D)
);

ninexnine_unit ninexnine_unit_4947(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2D00F),
				.b1(W2D01F),
				.b2(W2D02F),
				.b3(W2D10F),
				.b4(W2D11F),
				.b5(W2D12F),
				.b6(W2D20F),
				.b7(W2D21F),
				.b8(W2D22F),
				.c(c2F20D)
);

assign C220D=c2020D+c2120D+c2220D+c2320D+c2420D+c2520D+c2620D+c2720D+c2820D+c2920D+c2A20D+c2B20D+c2C20D+c2D20D+c2E20D+c2F20D;
assign A220D=(C220D>=0)?1:0;

assign P320D=A220D;

ninexnine_unit ninexnine_unit_4948(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2021D)
);

ninexnine_unit ninexnine_unit_4949(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2121D)
);

ninexnine_unit ninexnine_unit_4950(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2221D)
);

ninexnine_unit ninexnine_unit_4951(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2321D)
);

ninexnine_unit ninexnine_unit_4952(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2421D)
);

ninexnine_unit ninexnine_unit_4953(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2521D)
);

ninexnine_unit ninexnine_unit_4954(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2621D)
);

ninexnine_unit ninexnine_unit_4955(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2721D)
);

ninexnine_unit ninexnine_unit_4956(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2D008),
				.b1(W2D018),
				.b2(W2D028),
				.b3(W2D108),
				.b4(W2D118),
				.b5(W2D128),
				.b6(W2D208),
				.b7(W2D218),
				.b8(W2D228),
				.c(c2821D)
);

ninexnine_unit ninexnine_unit_4957(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2D009),
				.b1(W2D019),
				.b2(W2D029),
				.b3(W2D109),
				.b4(W2D119),
				.b5(W2D129),
				.b6(W2D209),
				.b7(W2D219),
				.b8(W2D229),
				.c(c2921D)
);

ninexnine_unit ninexnine_unit_4958(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2D00A),
				.b1(W2D01A),
				.b2(W2D02A),
				.b3(W2D10A),
				.b4(W2D11A),
				.b5(W2D12A),
				.b6(W2D20A),
				.b7(W2D21A),
				.b8(W2D22A),
				.c(c2A21D)
);

ninexnine_unit ninexnine_unit_4959(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2D00B),
				.b1(W2D01B),
				.b2(W2D02B),
				.b3(W2D10B),
				.b4(W2D11B),
				.b5(W2D12B),
				.b6(W2D20B),
				.b7(W2D21B),
				.b8(W2D22B),
				.c(c2B21D)
);

ninexnine_unit ninexnine_unit_4960(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2D00C),
				.b1(W2D01C),
				.b2(W2D02C),
				.b3(W2D10C),
				.b4(W2D11C),
				.b5(W2D12C),
				.b6(W2D20C),
				.b7(W2D21C),
				.b8(W2D22C),
				.c(c2C21D)
);

ninexnine_unit ninexnine_unit_4961(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2D00D),
				.b1(W2D01D),
				.b2(W2D02D),
				.b3(W2D10D),
				.b4(W2D11D),
				.b5(W2D12D),
				.b6(W2D20D),
				.b7(W2D21D),
				.b8(W2D22D),
				.c(c2D21D)
);

ninexnine_unit ninexnine_unit_4962(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2D00E),
				.b1(W2D01E),
				.b2(W2D02E),
				.b3(W2D10E),
				.b4(W2D11E),
				.b5(W2D12E),
				.b6(W2D20E),
				.b7(W2D21E),
				.b8(W2D22E),
				.c(c2E21D)
);

ninexnine_unit ninexnine_unit_4963(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2D00F),
				.b1(W2D01F),
				.b2(W2D02F),
				.b3(W2D10F),
				.b4(W2D11F),
				.b5(W2D12F),
				.b6(W2D20F),
				.b7(W2D21F),
				.b8(W2D22F),
				.c(c2F21D)
);

assign C221D=c2021D+c2121D+c2221D+c2321D+c2421D+c2521D+c2621D+c2721D+c2821D+c2921D+c2A21D+c2B21D+c2C21D+c2D21D+c2E21D+c2F21D;
assign A221D=(C221D>=0)?1:0;

assign P321D=A221D;

ninexnine_unit ninexnine_unit_4964(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2D000),
				.b1(W2D010),
				.b2(W2D020),
				.b3(W2D100),
				.b4(W2D110),
				.b5(W2D120),
				.b6(W2D200),
				.b7(W2D210),
				.b8(W2D220),
				.c(c2022D)
);

ninexnine_unit ninexnine_unit_4965(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2D001),
				.b1(W2D011),
				.b2(W2D021),
				.b3(W2D101),
				.b4(W2D111),
				.b5(W2D121),
				.b6(W2D201),
				.b7(W2D211),
				.b8(W2D221),
				.c(c2122D)
);

ninexnine_unit ninexnine_unit_4966(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2D002),
				.b1(W2D012),
				.b2(W2D022),
				.b3(W2D102),
				.b4(W2D112),
				.b5(W2D122),
				.b6(W2D202),
				.b7(W2D212),
				.b8(W2D222),
				.c(c2222D)
);

ninexnine_unit ninexnine_unit_4967(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2D003),
				.b1(W2D013),
				.b2(W2D023),
				.b3(W2D103),
				.b4(W2D113),
				.b5(W2D123),
				.b6(W2D203),
				.b7(W2D213),
				.b8(W2D223),
				.c(c2322D)
);

ninexnine_unit ninexnine_unit_4968(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2D004),
				.b1(W2D014),
				.b2(W2D024),
				.b3(W2D104),
				.b4(W2D114),
				.b5(W2D124),
				.b6(W2D204),
				.b7(W2D214),
				.b8(W2D224),
				.c(c2422D)
);

ninexnine_unit ninexnine_unit_4969(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2D005),
				.b1(W2D015),
				.b2(W2D025),
				.b3(W2D105),
				.b4(W2D115),
				.b5(W2D125),
				.b6(W2D205),
				.b7(W2D215),
				.b8(W2D225),
				.c(c2522D)
);

ninexnine_unit ninexnine_unit_4970(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2D006),
				.b1(W2D016),
				.b2(W2D026),
				.b3(W2D106),
				.b4(W2D116),
				.b5(W2D126),
				.b6(W2D206),
				.b7(W2D216),
				.b8(W2D226),
				.c(c2622D)
);

ninexnine_unit ninexnine_unit_4971(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2D007),
				.b1(W2D017),
				.b2(W2D027),
				.b3(W2D107),
				.b4(W2D117),
				.b5(W2D127),
				.b6(W2D207),
				.b7(W2D217),
				.b8(W2D227),
				.c(c2722D)
);

ninexnine_unit ninexnine_unit_4972(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2D008),
				.b1(W2D018),
				.b2(W2D028),
				.b3(W2D108),
				.b4(W2D118),
				.b5(W2D128),
				.b6(W2D208),
				.b7(W2D218),
				.b8(W2D228),
				.c(c2822D)
);

ninexnine_unit ninexnine_unit_4973(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2D009),
				.b1(W2D019),
				.b2(W2D029),
				.b3(W2D109),
				.b4(W2D119),
				.b5(W2D129),
				.b6(W2D209),
				.b7(W2D219),
				.b8(W2D229),
				.c(c2922D)
);

ninexnine_unit ninexnine_unit_4974(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2D00A),
				.b1(W2D01A),
				.b2(W2D02A),
				.b3(W2D10A),
				.b4(W2D11A),
				.b5(W2D12A),
				.b6(W2D20A),
				.b7(W2D21A),
				.b8(W2D22A),
				.c(c2A22D)
);

ninexnine_unit ninexnine_unit_4975(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2D00B),
				.b1(W2D01B),
				.b2(W2D02B),
				.b3(W2D10B),
				.b4(W2D11B),
				.b5(W2D12B),
				.b6(W2D20B),
				.b7(W2D21B),
				.b8(W2D22B),
				.c(c2B22D)
);

ninexnine_unit ninexnine_unit_4976(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2D00C),
				.b1(W2D01C),
				.b2(W2D02C),
				.b3(W2D10C),
				.b4(W2D11C),
				.b5(W2D12C),
				.b6(W2D20C),
				.b7(W2D21C),
				.b8(W2D22C),
				.c(c2C22D)
);

ninexnine_unit ninexnine_unit_4977(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2D00D),
				.b1(W2D01D),
				.b2(W2D02D),
				.b3(W2D10D),
				.b4(W2D11D),
				.b5(W2D12D),
				.b6(W2D20D),
				.b7(W2D21D),
				.b8(W2D22D),
				.c(c2D22D)
);

ninexnine_unit ninexnine_unit_4978(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2D00E),
				.b1(W2D01E),
				.b2(W2D02E),
				.b3(W2D10E),
				.b4(W2D11E),
				.b5(W2D12E),
				.b6(W2D20E),
				.b7(W2D21E),
				.b8(W2D22E),
				.c(c2E22D)
);

ninexnine_unit ninexnine_unit_4979(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2D00F),
				.b1(W2D01F),
				.b2(W2D02F),
				.b3(W2D10F),
				.b4(W2D11F),
				.b5(W2D12F),
				.b6(W2D20F),
				.b7(W2D21F),
				.b8(W2D22F),
				.c(c2F22D)
);

assign C222D=c2022D+c2122D+c2222D+c2322D+c2422D+c2522D+c2622D+c2722D+c2822D+c2922D+c2A22D+c2B22D+c2C22D+c2D22D+c2E22D+c2F22D;
assign A222D=(C222D>=0)?1:0;

assign P322D=A222D;

ninexnine_unit ninexnine_unit_4980(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2000E)
);

ninexnine_unit ninexnine_unit_4981(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2100E)
);

ninexnine_unit ninexnine_unit_4982(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2200E)
);

ninexnine_unit ninexnine_unit_4983(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2300E)
);

ninexnine_unit ninexnine_unit_4984(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2400E)
);

ninexnine_unit ninexnine_unit_4985(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2500E)
);

ninexnine_unit ninexnine_unit_4986(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2600E)
);

ninexnine_unit ninexnine_unit_4987(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2700E)
);

ninexnine_unit ninexnine_unit_4988(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2E008),
				.b1(W2E018),
				.b2(W2E028),
				.b3(W2E108),
				.b4(W2E118),
				.b5(W2E128),
				.b6(W2E208),
				.b7(W2E218),
				.b8(W2E228),
				.c(c2800E)
);

ninexnine_unit ninexnine_unit_4989(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2E009),
				.b1(W2E019),
				.b2(W2E029),
				.b3(W2E109),
				.b4(W2E119),
				.b5(W2E129),
				.b6(W2E209),
				.b7(W2E219),
				.b8(W2E229),
				.c(c2900E)
);

ninexnine_unit ninexnine_unit_4990(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2E00A),
				.b1(W2E01A),
				.b2(W2E02A),
				.b3(W2E10A),
				.b4(W2E11A),
				.b5(W2E12A),
				.b6(W2E20A),
				.b7(W2E21A),
				.b8(W2E22A),
				.c(c2A00E)
);

ninexnine_unit ninexnine_unit_4991(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2E00B),
				.b1(W2E01B),
				.b2(W2E02B),
				.b3(W2E10B),
				.b4(W2E11B),
				.b5(W2E12B),
				.b6(W2E20B),
				.b7(W2E21B),
				.b8(W2E22B),
				.c(c2B00E)
);

ninexnine_unit ninexnine_unit_4992(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2E00C),
				.b1(W2E01C),
				.b2(W2E02C),
				.b3(W2E10C),
				.b4(W2E11C),
				.b5(W2E12C),
				.b6(W2E20C),
				.b7(W2E21C),
				.b8(W2E22C),
				.c(c2C00E)
);

ninexnine_unit ninexnine_unit_4993(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2E00D),
				.b1(W2E01D),
				.b2(W2E02D),
				.b3(W2E10D),
				.b4(W2E11D),
				.b5(W2E12D),
				.b6(W2E20D),
				.b7(W2E21D),
				.b8(W2E22D),
				.c(c2D00E)
);

ninexnine_unit ninexnine_unit_4994(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2E00E),
				.b1(W2E01E),
				.b2(W2E02E),
				.b3(W2E10E),
				.b4(W2E11E),
				.b5(W2E12E),
				.b6(W2E20E),
				.b7(W2E21E),
				.b8(W2E22E),
				.c(c2E00E)
);

ninexnine_unit ninexnine_unit_4995(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2E00F),
				.b1(W2E01F),
				.b2(W2E02F),
				.b3(W2E10F),
				.b4(W2E11F),
				.b5(W2E12F),
				.b6(W2E20F),
				.b7(W2E21F),
				.b8(W2E22F),
				.c(c2F00E)
);

assign C200E=c2000E+c2100E+c2200E+c2300E+c2400E+c2500E+c2600E+c2700E+c2800E+c2900E+c2A00E+c2B00E+c2C00E+c2D00E+c2E00E+c2F00E;
assign A200E=(C200E>=0)?1:0;

assign P300E=A200E;

ninexnine_unit ninexnine_unit_4996(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2001E)
);

ninexnine_unit ninexnine_unit_4997(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2101E)
);

ninexnine_unit ninexnine_unit_4998(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2201E)
);

ninexnine_unit ninexnine_unit_4999(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2301E)
);

ninexnine_unit ninexnine_unit_5000(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2401E)
);

ninexnine_unit ninexnine_unit_5001(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2501E)
);

ninexnine_unit ninexnine_unit_5002(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2601E)
);

ninexnine_unit ninexnine_unit_5003(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2701E)
);

ninexnine_unit ninexnine_unit_5004(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2E008),
				.b1(W2E018),
				.b2(W2E028),
				.b3(W2E108),
				.b4(W2E118),
				.b5(W2E128),
				.b6(W2E208),
				.b7(W2E218),
				.b8(W2E228),
				.c(c2801E)
);

ninexnine_unit ninexnine_unit_5005(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2E009),
				.b1(W2E019),
				.b2(W2E029),
				.b3(W2E109),
				.b4(W2E119),
				.b5(W2E129),
				.b6(W2E209),
				.b7(W2E219),
				.b8(W2E229),
				.c(c2901E)
);

ninexnine_unit ninexnine_unit_5006(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2E00A),
				.b1(W2E01A),
				.b2(W2E02A),
				.b3(W2E10A),
				.b4(W2E11A),
				.b5(W2E12A),
				.b6(W2E20A),
				.b7(W2E21A),
				.b8(W2E22A),
				.c(c2A01E)
);

ninexnine_unit ninexnine_unit_5007(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2E00B),
				.b1(W2E01B),
				.b2(W2E02B),
				.b3(W2E10B),
				.b4(W2E11B),
				.b5(W2E12B),
				.b6(W2E20B),
				.b7(W2E21B),
				.b8(W2E22B),
				.c(c2B01E)
);

ninexnine_unit ninexnine_unit_5008(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2E00C),
				.b1(W2E01C),
				.b2(W2E02C),
				.b3(W2E10C),
				.b4(W2E11C),
				.b5(W2E12C),
				.b6(W2E20C),
				.b7(W2E21C),
				.b8(W2E22C),
				.c(c2C01E)
);

ninexnine_unit ninexnine_unit_5009(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2E00D),
				.b1(W2E01D),
				.b2(W2E02D),
				.b3(W2E10D),
				.b4(W2E11D),
				.b5(W2E12D),
				.b6(W2E20D),
				.b7(W2E21D),
				.b8(W2E22D),
				.c(c2D01E)
);

ninexnine_unit ninexnine_unit_5010(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2E00E),
				.b1(W2E01E),
				.b2(W2E02E),
				.b3(W2E10E),
				.b4(W2E11E),
				.b5(W2E12E),
				.b6(W2E20E),
				.b7(W2E21E),
				.b8(W2E22E),
				.c(c2E01E)
);

ninexnine_unit ninexnine_unit_5011(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2E00F),
				.b1(W2E01F),
				.b2(W2E02F),
				.b3(W2E10F),
				.b4(W2E11F),
				.b5(W2E12F),
				.b6(W2E20F),
				.b7(W2E21F),
				.b8(W2E22F),
				.c(c2F01E)
);

assign C201E=c2001E+c2101E+c2201E+c2301E+c2401E+c2501E+c2601E+c2701E+c2801E+c2901E+c2A01E+c2B01E+c2C01E+c2D01E+c2E01E+c2F01E;
assign A201E=(C201E>=0)?1:0;

assign P301E=A201E;

ninexnine_unit ninexnine_unit_5012(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2002E)
);

ninexnine_unit ninexnine_unit_5013(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2102E)
);

ninexnine_unit ninexnine_unit_5014(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2202E)
);

ninexnine_unit ninexnine_unit_5015(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2302E)
);

ninexnine_unit ninexnine_unit_5016(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2402E)
);

ninexnine_unit ninexnine_unit_5017(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2502E)
);

ninexnine_unit ninexnine_unit_5018(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2602E)
);

ninexnine_unit ninexnine_unit_5019(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2702E)
);

ninexnine_unit ninexnine_unit_5020(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2E008),
				.b1(W2E018),
				.b2(W2E028),
				.b3(W2E108),
				.b4(W2E118),
				.b5(W2E128),
				.b6(W2E208),
				.b7(W2E218),
				.b8(W2E228),
				.c(c2802E)
);

ninexnine_unit ninexnine_unit_5021(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2E009),
				.b1(W2E019),
				.b2(W2E029),
				.b3(W2E109),
				.b4(W2E119),
				.b5(W2E129),
				.b6(W2E209),
				.b7(W2E219),
				.b8(W2E229),
				.c(c2902E)
);

ninexnine_unit ninexnine_unit_5022(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2E00A),
				.b1(W2E01A),
				.b2(W2E02A),
				.b3(W2E10A),
				.b4(W2E11A),
				.b5(W2E12A),
				.b6(W2E20A),
				.b7(W2E21A),
				.b8(W2E22A),
				.c(c2A02E)
);

ninexnine_unit ninexnine_unit_5023(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2E00B),
				.b1(W2E01B),
				.b2(W2E02B),
				.b3(W2E10B),
				.b4(W2E11B),
				.b5(W2E12B),
				.b6(W2E20B),
				.b7(W2E21B),
				.b8(W2E22B),
				.c(c2B02E)
);

ninexnine_unit ninexnine_unit_5024(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2E00C),
				.b1(W2E01C),
				.b2(W2E02C),
				.b3(W2E10C),
				.b4(W2E11C),
				.b5(W2E12C),
				.b6(W2E20C),
				.b7(W2E21C),
				.b8(W2E22C),
				.c(c2C02E)
);

ninexnine_unit ninexnine_unit_5025(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2E00D),
				.b1(W2E01D),
				.b2(W2E02D),
				.b3(W2E10D),
				.b4(W2E11D),
				.b5(W2E12D),
				.b6(W2E20D),
				.b7(W2E21D),
				.b8(W2E22D),
				.c(c2D02E)
);

ninexnine_unit ninexnine_unit_5026(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2E00E),
				.b1(W2E01E),
				.b2(W2E02E),
				.b3(W2E10E),
				.b4(W2E11E),
				.b5(W2E12E),
				.b6(W2E20E),
				.b7(W2E21E),
				.b8(W2E22E),
				.c(c2E02E)
);

ninexnine_unit ninexnine_unit_5027(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2E00F),
				.b1(W2E01F),
				.b2(W2E02F),
				.b3(W2E10F),
				.b4(W2E11F),
				.b5(W2E12F),
				.b6(W2E20F),
				.b7(W2E21F),
				.b8(W2E22F),
				.c(c2F02E)
);

assign C202E=c2002E+c2102E+c2202E+c2302E+c2402E+c2502E+c2602E+c2702E+c2802E+c2902E+c2A02E+c2B02E+c2C02E+c2D02E+c2E02E+c2F02E;
assign A202E=(C202E>=0)?1:0;

assign P302E=A202E;

ninexnine_unit ninexnine_unit_5028(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2010E)
);

ninexnine_unit ninexnine_unit_5029(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2110E)
);

ninexnine_unit ninexnine_unit_5030(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2210E)
);

ninexnine_unit ninexnine_unit_5031(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2310E)
);

ninexnine_unit ninexnine_unit_5032(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2410E)
);

ninexnine_unit ninexnine_unit_5033(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2510E)
);

ninexnine_unit ninexnine_unit_5034(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2610E)
);

ninexnine_unit ninexnine_unit_5035(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2710E)
);

ninexnine_unit ninexnine_unit_5036(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2E008),
				.b1(W2E018),
				.b2(W2E028),
				.b3(W2E108),
				.b4(W2E118),
				.b5(W2E128),
				.b6(W2E208),
				.b7(W2E218),
				.b8(W2E228),
				.c(c2810E)
);

ninexnine_unit ninexnine_unit_5037(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2E009),
				.b1(W2E019),
				.b2(W2E029),
				.b3(W2E109),
				.b4(W2E119),
				.b5(W2E129),
				.b6(W2E209),
				.b7(W2E219),
				.b8(W2E229),
				.c(c2910E)
);

ninexnine_unit ninexnine_unit_5038(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2E00A),
				.b1(W2E01A),
				.b2(W2E02A),
				.b3(W2E10A),
				.b4(W2E11A),
				.b5(W2E12A),
				.b6(W2E20A),
				.b7(W2E21A),
				.b8(W2E22A),
				.c(c2A10E)
);

ninexnine_unit ninexnine_unit_5039(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2E00B),
				.b1(W2E01B),
				.b2(W2E02B),
				.b3(W2E10B),
				.b4(W2E11B),
				.b5(W2E12B),
				.b6(W2E20B),
				.b7(W2E21B),
				.b8(W2E22B),
				.c(c2B10E)
);

ninexnine_unit ninexnine_unit_5040(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2E00C),
				.b1(W2E01C),
				.b2(W2E02C),
				.b3(W2E10C),
				.b4(W2E11C),
				.b5(W2E12C),
				.b6(W2E20C),
				.b7(W2E21C),
				.b8(W2E22C),
				.c(c2C10E)
);

ninexnine_unit ninexnine_unit_5041(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2E00D),
				.b1(W2E01D),
				.b2(W2E02D),
				.b3(W2E10D),
				.b4(W2E11D),
				.b5(W2E12D),
				.b6(W2E20D),
				.b7(W2E21D),
				.b8(W2E22D),
				.c(c2D10E)
);

ninexnine_unit ninexnine_unit_5042(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2E00E),
				.b1(W2E01E),
				.b2(W2E02E),
				.b3(W2E10E),
				.b4(W2E11E),
				.b5(W2E12E),
				.b6(W2E20E),
				.b7(W2E21E),
				.b8(W2E22E),
				.c(c2E10E)
);

ninexnine_unit ninexnine_unit_5043(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2E00F),
				.b1(W2E01F),
				.b2(W2E02F),
				.b3(W2E10F),
				.b4(W2E11F),
				.b5(W2E12F),
				.b6(W2E20F),
				.b7(W2E21F),
				.b8(W2E22F),
				.c(c2F10E)
);

assign C210E=c2010E+c2110E+c2210E+c2310E+c2410E+c2510E+c2610E+c2710E+c2810E+c2910E+c2A10E+c2B10E+c2C10E+c2D10E+c2E10E+c2F10E;
assign A210E=(C210E>=0)?1:0;

assign P310E=A210E;

ninexnine_unit ninexnine_unit_5044(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2011E)
);

ninexnine_unit ninexnine_unit_5045(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2111E)
);

ninexnine_unit ninexnine_unit_5046(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2211E)
);

ninexnine_unit ninexnine_unit_5047(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2311E)
);

ninexnine_unit ninexnine_unit_5048(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2411E)
);

ninexnine_unit ninexnine_unit_5049(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2511E)
);

ninexnine_unit ninexnine_unit_5050(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2611E)
);

ninexnine_unit ninexnine_unit_5051(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2711E)
);

ninexnine_unit ninexnine_unit_5052(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2E008),
				.b1(W2E018),
				.b2(W2E028),
				.b3(W2E108),
				.b4(W2E118),
				.b5(W2E128),
				.b6(W2E208),
				.b7(W2E218),
				.b8(W2E228),
				.c(c2811E)
);

ninexnine_unit ninexnine_unit_5053(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2E009),
				.b1(W2E019),
				.b2(W2E029),
				.b3(W2E109),
				.b4(W2E119),
				.b5(W2E129),
				.b6(W2E209),
				.b7(W2E219),
				.b8(W2E229),
				.c(c2911E)
);

ninexnine_unit ninexnine_unit_5054(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2E00A),
				.b1(W2E01A),
				.b2(W2E02A),
				.b3(W2E10A),
				.b4(W2E11A),
				.b5(W2E12A),
				.b6(W2E20A),
				.b7(W2E21A),
				.b8(W2E22A),
				.c(c2A11E)
);

ninexnine_unit ninexnine_unit_5055(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2E00B),
				.b1(W2E01B),
				.b2(W2E02B),
				.b3(W2E10B),
				.b4(W2E11B),
				.b5(W2E12B),
				.b6(W2E20B),
				.b7(W2E21B),
				.b8(W2E22B),
				.c(c2B11E)
);

ninexnine_unit ninexnine_unit_5056(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2E00C),
				.b1(W2E01C),
				.b2(W2E02C),
				.b3(W2E10C),
				.b4(W2E11C),
				.b5(W2E12C),
				.b6(W2E20C),
				.b7(W2E21C),
				.b8(W2E22C),
				.c(c2C11E)
);

ninexnine_unit ninexnine_unit_5057(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2E00D),
				.b1(W2E01D),
				.b2(W2E02D),
				.b3(W2E10D),
				.b4(W2E11D),
				.b5(W2E12D),
				.b6(W2E20D),
				.b7(W2E21D),
				.b8(W2E22D),
				.c(c2D11E)
);

ninexnine_unit ninexnine_unit_5058(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2E00E),
				.b1(W2E01E),
				.b2(W2E02E),
				.b3(W2E10E),
				.b4(W2E11E),
				.b5(W2E12E),
				.b6(W2E20E),
				.b7(W2E21E),
				.b8(W2E22E),
				.c(c2E11E)
);

ninexnine_unit ninexnine_unit_5059(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2E00F),
				.b1(W2E01F),
				.b2(W2E02F),
				.b3(W2E10F),
				.b4(W2E11F),
				.b5(W2E12F),
				.b6(W2E20F),
				.b7(W2E21F),
				.b8(W2E22F),
				.c(c2F11E)
);

assign C211E=c2011E+c2111E+c2211E+c2311E+c2411E+c2511E+c2611E+c2711E+c2811E+c2911E+c2A11E+c2B11E+c2C11E+c2D11E+c2E11E+c2F11E;
assign A211E=(C211E>=0)?1:0;

assign P311E=A211E;

ninexnine_unit ninexnine_unit_5060(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2012E)
);

ninexnine_unit ninexnine_unit_5061(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2112E)
);

ninexnine_unit ninexnine_unit_5062(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2212E)
);

ninexnine_unit ninexnine_unit_5063(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2312E)
);

ninexnine_unit ninexnine_unit_5064(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2412E)
);

ninexnine_unit ninexnine_unit_5065(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2512E)
);

ninexnine_unit ninexnine_unit_5066(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2612E)
);

ninexnine_unit ninexnine_unit_5067(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2712E)
);

ninexnine_unit ninexnine_unit_5068(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2E008),
				.b1(W2E018),
				.b2(W2E028),
				.b3(W2E108),
				.b4(W2E118),
				.b5(W2E128),
				.b6(W2E208),
				.b7(W2E218),
				.b8(W2E228),
				.c(c2812E)
);

ninexnine_unit ninexnine_unit_5069(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2E009),
				.b1(W2E019),
				.b2(W2E029),
				.b3(W2E109),
				.b4(W2E119),
				.b5(W2E129),
				.b6(W2E209),
				.b7(W2E219),
				.b8(W2E229),
				.c(c2912E)
);

ninexnine_unit ninexnine_unit_5070(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2E00A),
				.b1(W2E01A),
				.b2(W2E02A),
				.b3(W2E10A),
				.b4(W2E11A),
				.b5(W2E12A),
				.b6(W2E20A),
				.b7(W2E21A),
				.b8(W2E22A),
				.c(c2A12E)
);

ninexnine_unit ninexnine_unit_5071(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2E00B),
				.b1(W2E01B),
				.b2(W2E02B),
				.b3(W2E10B),
				.b4(W2E11B),
				.b5(W2E12B),
				.b6(W2E20B),
				.b7(W2E21B),
				.b8(W2E22B),
				.c(c2B12E)
);

ninexnine_unit ninexnine_unit_5072(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2E00C),
				.b1(W2E01C),
				.b2(W2E02C),
				.b3(W2E10C),
				.b4(W2E11C),
				.b5(W2E12C),
				.b6(W2E20C),
				.b7(W2E21C),
				.b8(W2E22C),
				.c(c2C12E)
);

ninexnine_unit ninexnine_unit_5073(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2E00D),
				.b1(W2E01D),
				.b2(W2E02D),
				.b3(W2E10D),
				.b4(W2E11D),
				.b5(W2E12D),
				.b6(W2E20D),
				.b7(W2E21D),
				.b8(W2E22D),
				.c(c2D12E)
);

ninexnine_unit ninexnine_unit_5074(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2E00E),
				.b1(W2E01E),
				.b2(W2E02E),
				.b3(W2E10E),
				.b4(W2E11E),
				.b5(W2E12E),
				.b6(W2E20E),
				.b7(W2E21E),
				.b8(W2E22E),
				.c(c2E12E)
);

ninexnine_unit ninexnine_unit_5075(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2E00F),
				.b1(W2E01F),
				.b2(W2E02F),
				.b3(W2E10F),
				.b4(W2E11F),
				.b5(W2E12F),
				.b6(W2E20F),
				.b7(W2E21F),
				.b8(W2E22F),
				.c(c2F12E)
);

assign C212E=c2012E+c2112E+c2212E+c2312E+c2412E+c2512E+c2612E+c2712E+c2812E+c2912E+c2A12E+c2B12E+c2C12E+c2D12E+c2E12E+c2F12E;
assign A212E=(C212E>=0)?1:0;

assign P312E=A212E;

ninexnine_unit ninexnine_unit_5076(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2020E)
);

ninexnine_unit ninexnine_unit_5077(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2120E)
);

ninexnine_unit ninexnine_unit_5078(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2220E)
);

ninexnine_unit ninexnine_unit_5079(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2320E)
);

ninexnine_unit ninexnine_unit_5080(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2420E)
);

ninexnine_unit ninexnine_unit_5081(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2520E)
);

ninexnine_unit ninexnine_unit_5082(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2620E)
);

ninexnine_unit ninexnine_unit_5083(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2720E)
);

ninexnine_unit ninexnine_unit_5084(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2E008),
				.b1(W2E018),
				.b2(W2E028),
				.b3(W2E108),
				.b4(W2E118),
				.b5(W2E128),
				.b6(W2E208),
				.b7(W2E218),
				.b8(W2E228),
				.c(c2820E)
);

ninexnine_unit ninexnine_unit_5085(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2E009),
				.b1(W2E019),
				.b2(W2E029),
				.b3(W2E109),
				.b4(W2E119),
				.b5(W2E129),
				.b6(W2E209),
				.b7(W2E219),
				.b8(W2E229),
				.c(c2920E)
);

ninexnine_unit ninexnine_unit_5086(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2E00A),
				.b1(W2E01A),
				.b2(W2E02A),
				.b3(W2E10A),
				.b4(W2E11A),
				.b5(W2E12A),
				.b6(W2E20A),
				.b7(W2E21A),
				.b8(W2E22A),
				.c(c2A20E)
);

ninexnine_unit ninexnine_unit_5087(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2E00B),
				.b1(W2E01B),
				.b2(W2E02B),
				.b3(W2E10B),
				.b4(W2E11B),
				.b5(W2E12B),
				.b6(W2E20B),
				.b7(W2E21B),
				.b8(W2E22B),
				.c(c2B20E)
);

ninexnine_unit ninexnine_unit_5088(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2E00C),
				.b1(W2E01C),
				.b2(W2E02C),
				.b3(W2E10C),
				.b4(W2E11C),
				.b5(W2E12C),
				.b6(W2E20C),
				.b7(W2E21C),
				.b8(W2E22C),
				.c(c2C20E)
);

ninexnine_unit ninexnine_unit_5089(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2E00D),
				.b1(W2E01D),
				.b2(W2E02D),
				.b3(W2E10D),
				.b4(W2E11D),
				.b5(W2E12D),
				.b6(W2E20D),
				.b7(W2E21D),
				.b8(W2E22D),
				.c(c2D20E)
);

ninexnine_unit ninexnine_unit_5090(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2E00E),
				.b1(W2E01E),
				.b2(W2E02E),
				.b3(W2E10E),
				.b4(W2E11E),
				.b5(W2E12E),
				.b6(W2E20E),
				.b7(W2E21E),
				.b8(W2E22E),
				.c(c2E20E)
);

ninexnine_unit ninexnine_unit_5091(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2E00F),
				.b1(W2E01F),
				.b2(W2E02F),
				.b3(W2E10F),
				.b4(W2E11F),
				.b5(W2E12F),
				.b6(W2E20F),
				.b7(W2E21F),
				.b8(W2E22F),
				.c(c2F20E)
);

assign C220E=c2020E+c2120E+c2220E+c2320E+c2420E+c2520E+c2620E+c2720E+c2820E+c2920E+c2A20E+c2B20E+c2C20E+c2D20E+c2E20E+c2F20E;
assign A220E=(C220E>=0)?1:0;

assign P320E=A220E;

ninexnine_unit ninexnine_unit_5092(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2021E)
);

ninexnine_unit ninexnine_unit_5093(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2121E)
);

ninexnine_unit ninexnine_unit_5094(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2221E)
);

ninexnine_unit ninexnine_unit_5095(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2321E)
);

ninexnine_unit ninexnine_unit_5096(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2421E)
);

ninexnine_unit ninexnine_unit_5097(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2521E)
);

ninexnine_unit ninexnine_unit_5098(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2621E)
);

ninexnine_unit ninexnine_unit_5099(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2721E)
);

ninexnine_unit ninexnine_unit_5100(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2E008),
				.b1(W2E018),
				.b2(W2E028),
				.b3(W2E108),
				.b4(W2E118),
				.b5(W2E128),
				.b6(W2E208),
				.b7(W2E218),
				.b8(W2E228),
				.c(c2821E)
);

ninexnine_unit ninexnine_unit_5101(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2E009),
				.b1(W2E019),
				.b2(W2E029),
				.b3(W2E109),
				.b4(W2E119),
				.b5(W2E129),
				.b6(W2E209),
				.b7(W2E219),
				.b8(W2E229),
				.c(c2921E)
);

ninexnine_unit ninexnine_unit_5102(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2E00A),
				.b1(W2E01A),
				.b2(W2E02A),
				.b3(W2E10A),
				.b4(W2E11A),
				.b5(W2E12A),
				.b6(W2E20A),
				.b7(W2E21A),
				.b8(W2E22A),
				.c(c2A21E)
);

ninexnine_unit ninexnine_unit_5103(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2E00B),
				.b1(W2E01B),
				.b2(W2E02B),
				.b3(W2E10B),
				.b4(W2E11B),
				.b5(W2E12B),
				.b6(W2E20B),
				.b7(W2E21B),
				.b8(W2E22B),
				.c(c2B21E)
);

ninexnine_unit ninexnine_unit_5104(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2E00C),
				.b1(W2E01C),
				.b2(W2E02C),
				.b3(W2E10C),
				.b4(W2E11C),
				.b5(W2E12C),
				.b6(W2E20C),
				.b7(W2E21C),
				.b8(W2E22C),
				.c(c2C21E)
);

ninexnine_unit ninexnine_unit_5105(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2E00D),
				.b1(W2E01D),
				.b2(W2E02D),
				.b3(W2E10D),
				.b4(W2E11D),
				.b5(W2E12D),
				.b6(W2E20D),
				.b7(W2E21D),
				.b8(W2E22D),
				.c(c2D21E)
);

ninexnine_unit ninexnine_unit_5106(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2E00E),
				.b1(W2E01E),
				.b2(W2E02E),
				.b3(W2E10E),
				.b4(W2E11E),
				.b5(W2E12E),
				.b6(W2E20E),
				.b7(W2E21E),
				.b8(W2E22E),
				.c(c2E21E)
);

ninexnine_unit ninexnine_unit_5107(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2E00F),
				.b1(W2E01F),
				.b2(W2E02F),
				.b3(W2E10F),
				.b4(W2E11F),
				.b5(W2E12F),
				.b6(W2E20F),
				.b7(W2E21F),
				.b8(W2E22F),
				.c(c2F21E)
);

assign C221E=c2021E+c2121E+c2221E+c2321E+c2421E+c2521E+c2621E+c2721E+c2821E+c2921E+c2A21E+c2B21E+c2C21E+c2D21E+c2E21E+c2F21E;
assign A221E=(C221E>=0)?1:0;

assign P321E=A221E;

ninexnine_unit ninexnine_unit_5108(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2E000),
				.b1(W2E010),
				.b2(W2E020),
				.b3(W2E100),
				.b4(W2E110),
				.b5(W2E120),
				.b6(W2E200),
				.b7(W2E210),
				.b8(W2E220),
				.c(c2022E)
);

ninexnine_unit ninexnine_unit_5109(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2E001),
				.b1(W2E011),
				.b2(W2E021),
				.b3(W2E101),
				.b4(W2E111),
				.b5(W2E121),
				.b6(W2E201),
				.b7(W2E211),
				.b8(W2E221),
				.c(c2122E)
);

ninexnine_unit ninexnine_unit_5110(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2E002),
				.b1(W2E012),
				.b2(W2E022),
				.b3(W2E102),
				.b4(W2E112),
				.b5(W2E122),
				.b6(W2E202),
				.b7(W2E212),
				.b8(W2E222),
				.c(c2222E)
);

ninexnine_unit ninexnine_unit_5111(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2E003),
				.b1(W2E013),
				.b2(W2E023),
				.b3(W2E103),
				.b4(W2E113),
				.b5(W2E123),
				.b6(W2E203),
				.b7(W2E213),
				.b8(W2E223),
				.c(c2322E)
);

ninexnine_unit ninexnine_unit_5112(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2E004),
				.b1(W2E014),
				.b2(W2E024),
				.b3(W2E104),
				.b4(W2E114),
				.b5(W2E124),
				.b6(W2E204),
				.b7(W2E214),
				.b8(W2E224),
				.c(c2422E)
);

ninexnine_unit ninexnine_unit_5113(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2E005),
				.b1(W2E015),
				.b2(W2E025),
				.b3(W2E105),
				.b4(W2E115),
				.b5(W2E125),
				.b6(W2E205),
				.b7(W2E215),
				.b8(W2E225),
				.c(c2522E)
);

ninexnine_unit ninexnine_unit_5114(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2E006),
				.b1(W2E016),
				.b2(W2E026),
				.b3(W2E106),
				.b4(W2E116),
				.b5(W2E126),
				.b6(W2E206),
				.b7(W2E216),
				.b8(W2E226),
				.c(c2622E)
);

ninexnine_unit ninexnine_unit_5115(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2E007),
				.b1(W2E017),
				.b2(W2E027),
				.b3(W2E107),
				.b4(W2E117),
				.b5(W2E127),
				.b6(W2E207),
				.b7(W2E217),
				.b8(W2E227),
				.c(c2722E)
);

ninexnine_unit ninexnine_unit_5116(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2E008),
				.b1(W2E018),
				.b2(W2E028),
				.b3(W2E108),
				.b4(W2E118),
				.b5(W2E128),
				.b6(W2E208),
				.b7(W2E218),
				.b8(W2E228),
				.c(c2822E)
);

ninexnine_unit ninexnine_unit_5117(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2E009),
				.b1(W2E019),
				.b2(W2E029),
				.b3(W2E109),
				.b4(W2E119),
				.b5(W2E129),
				.b6(W2E209),
				.b7(W2E219),
				.b8(W2E229),
				.c(c2922E)
);

ninexnine_unit ninexnine_unit_5118(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2E00A),
				.b1(W2E01A),
				.b2(W2E02A),
				.b3(W2E10A),
				.b4(W2E11A),
				.b5(W2E12A),
				.b6(W2E20A),
				.b7(W2E21A),
				.b8(W2E22A),
				.c(c2A22E)
);

ninexnine_unit ninexnine_unit_5119(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2E00B),
				.b1(W2E01B),
				.b2(W2E02B),
				.b3(W2E10B),
				.b4(W2E11B),
				.b5(W2E12B),
				.b6(W2E20B),
				.b7(W2E21B),
				.b8(W2E22B),
				.c(c2B22E)
);

ninexnine_unit ninexnine_unit_5120(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2E00C),
				.b1(W2E01C),
				.b2(W2E02C),
				.b3(W2E10C),
				.b4(W2E11C),
				.b5(W2E12C),
				.b6(W2E20C),
				.b7(W2E21C),
				.b8(W2E22C),
				.c(c2C22E)
);

ninexnine_unit ninexnine_unit_5121(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2E00D),
				.b1(W2E01D),
				.b2(W2E02D),
				.b3(W2E10D),
				.b4(W2E11D),
				.b5(W2E12D),
				.b6(W2E20D),
				.b7(W2E21D),
				.b8(W2E22D),
				.c(c2D22E)
);

ninexnine_unit ninexnine_unit_5122(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2E00E),
				.b1(W2E01E),
				.b2(W2E02E),
				.b3(W2E10E),
				.b4(W2E11E),
				.b5(W2E12E),
				.b6(W2E20E),
				.b7(W2E21E),
				.b8(W2E22E),
				.c(c2E22E)
);

ninexnine_unit ninexnine_unit_5123(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2E00F),
				.b1(W2E01F),
				.b2(W2E02F),
				.b3(W2E10F),
				.b4(W2E11F),
				.b5(W2E12F),
				.b6(W2E20F),
				.b7(W2E21F),
				.b8(W2E22F),
				.c(c2F22E)
);

assign C222E=c2022E+c2122E+c2222E+c2322E+c2422E+c2522E+c2622E+c2722E+c2822E+c2922E+c2A22E+c2B22E+c2C22E+c2D22E+c2E22E+c2F22E;
assign A222E=(C222E>=0)?1:0;

assign P322E=A222E;

ninexnine_unit ninexnine_unit_5124(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2000F)
);

ninexnine_unit ninexnine_unit_5125(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2100F)
);

ninexnine_unit ninexnine_unit_5126(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2200F)
);

ninexnine_unit ninexnine_unit_5127(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2300F)
);

ninexnine_unit ninexnine_unit_5128(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2400F)
);

ninexnine_unit ninexnine_unit_5129(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2500F)
);

ninexnine_unit ninexnine_unit_5130(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2600F)
);

ninexnine_unit ninexnine_unit_5131(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2700F)
);

ninexnine_unit ninexnine_unit_5132(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2F008),
				.b1(W2F018),
				.b2(W2F028),
				.b3(W2F108),
				.b4(W2F118),
				.b5(W2F128),
				.b6(W2F208),
				.b7(W2F218),
				.b8(W2F228),
				.c(c2800F)
);

ninexnine_unit ninexnine_unit_5133(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2F009),
				.b1(W2F019),
				.b2(W2F029),
				.b3(W2F109),
				.b4(W2F119),
				.b5(W2F129),
				.b6(W2F209),
				.b7(W2F219),
				.b8(W2F229),
				.c(c2900F)
);

ninexnine_unit ninexnine_unit_5134(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2F00A),
				.b1(W2F01A),
				.b2(W2F02A),
				.b3(W2F10A),
				.b4(W2F11A),
				.b5(W2F12A),
				.b6(W2F20A),
				.b7(W2F21A),
				.b8(W2F22A),
				.c(c2A00F)
);

ninexnine_unit ninexnine_unit_5135(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2F00B),
				.b1(W2F01B),
				.b2(W2F02B),
				.b3(W2F10B),
				.b4(W2F11B),
				.b5(W2F12B),
				.b6(W2F20B),
				.b7(W2F21B),
				.b8(W2F22B),
				.c(c2B00F)
);

ninexnine_unit ninexnine_unit_5136(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2F00C),
				.b1(W2F01C),
				.b2(W2F02C),
				.b3(W2F10C),
				.b4(W2F11C),
				.b5(W2F12C),
				.b6(W2F20C),
				.b7(W2F21C),
				.b8(W2F22C),
				.c(c2C00F)
);

ninexnine_unit ninexnine_unit_5137(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2F00D),
				.b1(W2F01D),
				.b2(W2F02D),
				.b3(W2F10D),
				.b4(W2F11D),
				.b5(W2F12D),
				.b6(W2F20D),
				.b7(W2F21D),
				.b8(W2F22D),
				.c(c2D00F)
);

ninexnine_unit ninexnine_unit_5138(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2F00E),
				.b1(W2F01E),
				.b2(W2F02E),
				.b3(W2F10E),
				.b4(W2F11E),
				.b5(W2F12E),
				.b6(W2F20E),
				.b7(W2F21E),
				.b8(W2F22E),
				.c(c2E00F)
);

ninexnine_unit ninexnine_unit_5139(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2F00F),
				.b1(W2F01F),
				.b2(W2F02F),
				.b3(W2F10F),
				.b4(W2F11F),
				.b5(W2F12F),
				.b6(W2F20F),
				.b7(W2F21F),
				.b8(W2F22F),
				.c(c2F00F)
);

assign C200F=c2000F+c2100F+c2200F+c2300F+c2400F+c2500F+c2600F+c2700F+c2800F+c2900F+c2A00F+c2B00F+c2C00F+c2D00F+c2E00F+c2F00F;
assign A200F=(C200F>=0)?1:0;

assign P300F=A200F;

ninexnine_unit ninexnine_unit_5140(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2001F)
);

ninexnine_unit ninexnine_unit_5141(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2101F)
);

ninexnine_unit ninexnine_unit_5142(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2201F)
);

ninexnine_unit ninexnine_unit_5143(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2301F)
);

ninexnine_unit ninexnine_unit_5144(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2401F)
);

ninexnine_unit ninexnine_unit_5145(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2501F)
);

ninexnine_unit ninexnine_unit_5146(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2601F)
);

ninexnine_unit ninexnine_unit_5147(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2701F)
);

ninexnine_unit ninexnine_unit_5148(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2F008),
				.b1(W2F018),
				.b2(W2F028),
				.b3(W2F108),
				.b4(W2F118),
				.b5(W2F128),
				.b6(W2F208),
				.b7(W2F218),
				.b8(W2F228),
				.c(c2801F)
);

ninexnine_unit ninexnine_unit_5149(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2F009),
				.b1(W2F019),
				.b2(W2F029),
				.b3(W2F109),
				.b4(W2F119),
				.b5(W2F129),
				.b6(W2F209),
				.b7(W2F219),
				.b8(W2F229),
				.c(c2901F)
);

ninexnine_unit ninexnine_unit_5150(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2F00A),
				.b1(W2F01A),
				.b2(W2F02A),
				.b3(W2F10A),
				.b4(W2F11A),
				.b5(W2F12A),
				.b6(W2F20A),
				.b7(W2F21A),
				.b8(W2F22A),
				.c(c2A01F)
);

ninexnine_unit ninexnine_unit_5151(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2F00B),
				.b1(W2F01B),
				.b2(W2F02B),
				.b3(W2F10B),
				.b4(W2F11B),
				.b5(W2F12B),
				.b6(W2F20B),
				.b7(W2F21B),
				.b8(W2F22B),
				.c(c2B01F)
);

ninexnine_unit ninexnine_unit_5152(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2F00C),
				.b1(W2F01C),
				.b2(W2F02C),
				.b3(W2F10C),
				.b4(W2F11C),
				.b5(W2F12C),
				.b6(W2F20C),
				.b7(W2F21C),
				.b8(W2F22C),
				.c(c2C01F)
);

ninexnine_unit ninexnine_unit_5153(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2F00D),
				.b1(W2F01D),
				.b2(W2F02D),
				.b3(W2F10D),
				.b4(W2F11D),
				.b5(W2F12D),
				.b6(W2F20D),
				.b7(W2F21D),
				.b8(W2F22D),
				.c(c2D01F)
);

ninexnine_unit ninexnine_unit_5154(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2F00E),
				.b1(W2F01E),
				.b2(W2F02E),
				.b3(W2F10E),
				.b4(W2F11E),
				.b5(W2F12E),
				.b6(W2F20E),
				.b7(W2F21E),
				.b8(W2F22E),
				.c(c2E01F)
);

ninexnine_unit ninexnine_unit_5155(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2F00F),
				.b1(W2F01F),
				.b2(W2F02F),
				.b3(W2F10F),
				.b4(W2F11F),
				.b5(W2F12F),
				.b6(W2F20F),
				.b7(W2F21F),
				.b8(W2F22F),
				.c(c2F01F)
);

assign C201F=c2001F+c2101F+c2201F+c2301F+c2401F+c2501F+c2601F+c2701F+c2801F+c2901F+c2A01F+c2B01F+c2C01F+c2D01F+c2E01F+c2F01F;
assign A201F=(C201F>=0)?1:0;

assign P301F=A201F;

ninexnine_unit ninexnine_unit_5156(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2002F)
);

ninexnine_unit ninexnine_unit_5157(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2102F)
);

ninexnine_unit ninexnine_unit_5158(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2202F)
);

ninexnine_unit ninexnine_unit_5159(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2302F)
);

ninexnine_unit ninexnine_unit_5160(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2402F)
);

ninexnine_unit ninexnine_unit_5161(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2502F)
);

ninexnine_unit ninexnine_unit_5162(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2602F)
);

ninexnine_unit ninexnine_unit_5163(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2702F)
);

ninexnine_unit ninexnine_unit_5164(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2F008),
				.b1(W2F018),
				.b2(W2F028),
				.b3(W2F108),
				.b4(W2F118),
				.b5(W2F128),
				.b6(W2F208),
				.b7(W2F218),
				.b8(W2F228),
				.c(c2802F)
);

ninexnine_unit ninexnine_unit_5165(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2F009),
				.b1(W2F019),
				.b2(W2F029),
				.b3(W2F109),
				.b4(W2F119),
				.b5(W2F129),
				.b6(W2F209),
				.b7(W2F219),
				.b8(W2F229),
				.c(c2902F)
);

ninexnine_unit ninexnine_unit_5166(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2F00A),
				.b1(W2F01A),
				.b2(W2F02A),
				.b3(W2F10A),
				.b4(W2F11A),
				.b5(W2F12A),
				.b6(W2F20A),
				.b7(W2F21A),
				.b8(W2F22A),
				.c(c2A02F)
);

ninexnine_unit ninexnine_unit_5167(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2F00B),
				.b1(W2F01B),
				.b2(W2F02B),
				.b3(W2F10B),
				.b4(W2F11B),
				.b5(W2F12B),
				.b6(W2F20B),
				.b7(W2F21B),
				.b8(W2F22B),
				.c(c2B02F)
);

ninexnine_unit ninexnine_unit_5168(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2F00C),
				.b1(W2F01C),
				.b2(W2F02C),
				.b3(W2F10C),
				.b4(W2F11C),
				.b5(W2F12C),
				.b6(W2F20C),
				.b7(W2F21C),
				.b8(W2F22C),
				.c(c2C02F)
);

ninexnine_unit ninexnine_unit_5169(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2F00D),
				.b1(W2F01D),
				.b2(W2F02D),
				.b3(W2F10D),
				.b4(W2F11D),
				.b5(W2F12D),
				.b6(W2F20D),
				.b7(W2F21D),
				.b8(W2F22D),
				.c(c2D02F)
);

ninexnine_unit ninexnine_unit_5170(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2F00E),
				.b1(W2F01E),
				.b2(W2F02E),
				.b3(W2F10E),
				.b4(W2F11E),
				.b5(W2F12E),
				.b6(W2F20E),
				.b7(W2F21E),
				.b8(W2F22E),
				.c(c2E02F)
);

ninexnine_unit ninexnine_unit_5171(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2F00F),
				.b1(W2F01F),
				.b2(W2F02F),
				.b3(W2F10F),
				.b4(W2F11F),
				.b5(W2F12F),
				.b6(W2F20F),
				.b7(W2F21F),
				.b8(W2F22F),
				.c(c2F02F)
);

assign C202F=c2002F+c2102F+c2202F+c2302F+c2402F+c2502F+c2602F+c2702F+c2802F+c2902F+c2A02F+c2B02F+c2C02F+c2D02F+c2E02F+c2F02F;
assign A202F=(C202F>=0)?1:0;

assign P302F=A202F;

ninexnine_unit ninexnine_unit_5172(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2010F)
);

ninexnine_unit ninexnine_unit_5173(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2110F)
);

ninexnine_unit ninexnine_unit_5174(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2210F)
);

ninexnine_unit ninexnine_unit_5175(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2310F)
);

ninexnine_unit ninexnine_unit_5176(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2410F)
);

ninexnine_unit ninexnine_unit_5177(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2510F)
);

ninexnine_unit ninexnine_unit_5178(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2610F)
);

ninexnine_unit ninexnine_unit_5179(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2710F)
);

ninexnine_unit ninexnine_unit_5180(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2F008),
				.b1(W2F018),
				.b2(W2F028),
				.b3(W2F108),
				.b4(W2F118),
				.b5(W2F128),
				.b6(W2F208),
				.b7(W2F218),
				.b8(W2F228),
				.c(c2810F)
);

ninexnine_unit ninexnine_unit_5181(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2F009),
				.b1(W2F019),
				.b2(W2F029),
				.b3(W2F109),
				.b4(W2F119),
				.b5(W2F129),
				.b6(W2F209),
				.b7(W2F219),
				.b8(W2F229),
				.c(c2910F)
);

ninexnine_unit ninexnine_unit_5182(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2F00A),
				.b1(W2F01A),
				.b2(W2F02A),
				.b3(W2F10A),
				.b4(W2F11A),
				.b5(W2F12A),
				.b6(W2F20A),
				.b7(W2F21A),
				.b8(W2F22A),
				.c(c2A10F)
);

ninexnine_unit ninexnine_unit_5183(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2F00B),
				.b1(W2F01B),
				.b2(W2F02B),
				.b3(W2F10B),
				.b4(W2F11B),
				.b5(W2F12B),
				.b6(W2F20B),
				.b7(W2F21B),
				.b8(W2F22B),
				.c(c2B10F)
);

ninexnine_unit ninexnine_unit_5184(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2F00C),
				.b1(W2F01C),
				.b2(W2F02C),
				.b3(W2F10C),
				.b4(W2F11C),
				.b5(W2F12C),
				.b6(W2F20C),
				.b7(W2F21C),
				.b8(W2F22C),
				.c(c2C10F)
);

ninexnine_unit ninexnine_unit_5185(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2F00D),
				.b1(W2F01D),
				.b2(W2F02D),
				.b3(W2F10D),
				.b4(W2F11D),
				.b5(W2F12D),
				.b6(W2F20D),
				.b7(W2F21D),
				.b8(W2F22D),
				.c(c2D10F)
);

ninexnine_unit ninexnine_unit_5186(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2F00E),
				.b1(W2F01E),
				.b2(W2F02E),
				.b3(W2F10E),
				.b4(W2F11E),
				.b5(W2F12E),
				.b6(W2F20E),
				.b7(W2F21E),
				.b8(W2F22E),
				.c(c2E10F)
);

ninexnine_unit ninexnine_unit_5187(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2F00F),
				.b1(W2F01F),
				.b2(W2F02F),
				.b3(W2F10F),
				.b4(W2F11F),
				.b5(W2F12F),
				.b6(W2F20F),
				.b7(W2F21F),
				.b8(W2F22F),
				.c(c2F10F)
);

assign C210F=c2010F+c2110F+c2210F+c2310F+c2410F+c2510F+c2610F+c2710F+c2810F+c2910F+c2A10F+c2B10F+c2C10F+c2D10F+c2E10F+c2F10F;
assign A210F=(C210F>=0)?1:0;

assign P310F=A210F;

ninexnine_unit ninexnine_unit_5188(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2011F)
);

ninexnine_unit ninexnine_unit_5189(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2111F)
);

ninexnine_unit ninexnine_unit_5190(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2211F)
);

ninexnine_unit ninexnine_unit_5191(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2311F)
);

ninexnine_unit ninexnine_unit_5192(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2411F)
);

ninexnine_unit ninexnine_unit_5193(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2511F)
);

ninexnine_unit ninexnine_unit_5194(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2611F)
);

ninexnine_unit ninexnine_unit_5195(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2711F)
);

ninexnine_unit ninexnine_unit_5196(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2F008),
				.b1(W2F018),
				.b2(W2F028),
				.b3(W2F108),
				.b4(W2F118),
				.b5(W2F128),
				.b6(W2F208),
				.b7(W2F218),
				.b8(W2F228),
				.c(c2811F)
);

ninexnine_unit ninexnine_unit_5197(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2F009),
				.b1(W2F019),
				.b2(W2F029),
				.b3(W2F109),
				.b4(W2F119),
				.b5(W2F129),
				.b6(W2F209),
				.b7(W2F219),
				.b8(W2F229),
				.c(c2911F)
);

ninexnine_unit ninexnine_unit_5198(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2F00A),
				.b1(W2F01A),
				.b2(W2F02A),
				.b3(W2F10A),
				.b4(W2F11A),
				.b5(W2F12A),
				.b6(W2F20A),
				.b7(W2F21A),
				.b8(W2F22A),
				.c(c2A11F)
);

ninexnine_unit ninexnine_unit_5199(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2F00B),
				.b1(W2F01B),
				.b2(W2F02B),
				.b3(W2F10B),
				.b4(W2F11B),
				.b5(W2F12B),
				.b6(W2F20B),
				.b7(W2F21B),
				.b8(W2F22B),
				.c(c2B11F)
);

ninexnine_unit ninexnine_unit_5200(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2F00C),
				.b1(W2F01C),
				.b2(W2F02C),
				.b3(W2F10C),
				.b4(W2F11C),
				.b5(W2F12C),
				.b6(W2F20C),
				.b7(W2F21C),
				.b8(W2F22C),
				.c(c2C11F)
);

ninexnine_unit ninexnine_unit_5201(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2F00D),
				.b1(W2F01D),
				.b2(W2F02D),
				.b3(W2F10D),
				.b4(W2F11D),
				.b5(W2F12D),
				.b6(W2F20D),
				.b7(W2F21D),
				.b8(W2F22D),
				.c(c2D11F)
);

ninexnine_unit ninexnine_unit_5202(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2F00E),
				.b1(W2F01E),
				.b2(W2F02E),
				.b3(W2F10E),
				.b4(W2F11E),
				.b5(W2F12E),
				.b6(W2F20E),
				.b7(W2F21E),
				.b8(W2F22E),
				.c(c2E11F)
);

ninexnine_unit ninexnine_unit_5203(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2F00F),
				.b1(W2F01F),
				.b2(W2F02F),
				.b3(W2F10F),
				.b4(W2F11F),
				.b5(W2F12F),
				.b6(W2F20F),
				.b7(W2F21F),
				.b8(W2F22F),
				.c(c2F11F)
);

assign C211F=c2011F+c2111F+c2211F+c2311F+c2411F+c2511F+c2611F+c2711F+c2811F+c2911F+c2A11F+c2B11F+c2C11F+c2D11F+c2E11F+c2F11F;
assign A211F=(C211F>=0)?1:0;

assign P311F=A211F;

ninexnine_unit ninexnine_unit_5204(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2012F)
);

ninexnine_unit ninexnine_unit_5205(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2112F)
);

ninexnine_unit ninexnine_unit_5206(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2212F)
);

ninexnine_unit ninexnine_unit_5207(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2312F)
);

ninexnine_unit ninexnine_unit_5208(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2412F)
);

ninexnine_unit ninexnine_unit_5209(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2512F)
);

ninexnine_unit ninexnine_unit_5210(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2612F)
);

ninexnine_unit ninexnine_unit_5211(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2712F)
);

ninexnine_unit ninexnine_unit_5212(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2F008),
				.b1(W2F018),
				.b2(W2F028),
				.b3(W2F108),
				.b4(W2F118),
				.b5(W2F128),
				.b6(W2F208),
				.b7(W2F218),
				.b8(W2F228),
				.c(c2812F)
);

ninexnine_unit ninexnine_unit_5213(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2F009),
				.b1(W2F019),
				.b2(W2F029),
				.b3(W2F109),
				.b4(W2F119),
				.b5(W2F129),
				.b6(W2F209),
				.b7(W2F219),
				.b8(W2F229),
				.c(c2912F)
);

ninexnine_unit ninexnine_unit_5214(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2F00A),
				.b1(W2F01A),
				.b2(W2F02A),
				.b3(W2F10A),
				.b4(W2F11A),
				.b5(W2F12A),
				.b6(W2F20A),
				.b7(W2F21A),
				.b8(W2F22A),
				.c(c2A12F)
);

ninexnine_unit ninexnine_unit_5215(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2F00B),
				.b1(W2F01B),
				.b2(W2F02B),
				.b3(W2F10B),
				.b4(W2F11B),
				.b5(W2F12B),
				.b6(W2F20B),
				.b7(W2F21B),
				.b8(W2F22B),
				.c(c2B12F)
);

ninexnine_unit ninexnine_unit_5216(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2F00C),
				.b1(W2F01C),
				.b2(W2F02C),
				.b3(W2F10C),
				.b4(W2F11C),
				.b5(W2F12C),
				.b6(W2F20C),
				.b7(W2F21C),
				.b8(W2F22C),
				.c(c2C12F)
);

ninexnine_unit ninexnine_unit_5217(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2F00D),
				.b1(W2F01D),
				.b2(W2F02D),
				.b3(W2F10D),
				.b4(W2F11D),
				.b5(W2F12D),
				.b6(W2F20D),
				.b7(W2F21D),
				.b8(W2F22D),
				.c(c2D12F)
);

ninexnine_unit ninexnine_unit_5218(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2F00E),
				.b1(W2F01E),
				.b2(W2F02E),
				.b3(W2F10E),
				.b4(W2F11E),
				.b5(W2F12E),
				.b6(W2F20E),
				.b7(W2F21E),
				.b8(W2F22E),
				.c(c2E12F)
);

ninexnine_unit ninexnine_unit_5219(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2F00F),
				.b1(W2F01F),
				.b2(W2F02F),
				.b3(W2F10F),
				.b4(W2F11F),
				.b5(W2F12F),
				.b6(W2F20F),
				.b7(W2F21F),
				.b8(W2F22F),
				.c(c2F12F)
);

assign C212F=c2012F+c2112F+c2212F+c2312F+c2412F+c2512F+c2612F+c2712F+c2812F+c2912F+c2A12F+c2B12F+c2C12F+c2D12F+c2E12F+c2F12F;
assign A212F=(C212F>=0)?1:0;

assign P312F=A212F;

ninexnine_unit ninexnine_unit_5220(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2020F)
);

ninexnine_unit ninexnine_unit_5221(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2120F)
);

ninexnine_unit ninexnine_unit_5222(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2220F)
);

ninexnine_unit ninexnine_unit_5223(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2320F)
);

ninexnine_unit ninexnine_unit_5224(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2420F)
);

ninexnine_unit ninexnine_unit_5225(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2520F)
);

ninexnine_unit ninexnine_unit_5226(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2620F)
);

ninexnine_unit ninexnine_unit_5227(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2720F)
);

ninexnine_unit ninexnine_unit_5228(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2F008),
				.b1(W2F018),
				.b2(W2F028),
				.b3(W2F108),
				.b4(W2F118),
				.b5(W2F128),
				.b6(W2F208),
				.b7(W2F218),
				.b8(W2F228),
				.c(c2820F)
);

ninexnine_unit ninexnine_unit_5229(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2F009),
				.b1(W2F019),
				.b2(W2F029),
				.b3(W2F109),
				.b4(W2F119),
				.b5(W2F129),
				.b6(W2F209),
				.b7(W2F219),
				.b8(W2F229),
				.c(c2920F)
);

ninexnine_unit ninexnine_unit_5230(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2F00A),
				.b1(W2F01A),
				.b2(W2F02A),
				.b3(W2F10A),
				.b4(W2F11A),
				.b5(W2F12A),
				.b6(W2F20A),
				.b7(W2F21A),
				.b8(W2F22A),
				.c(c2A20F)
);

ninexnine_unit ninexnine_unit_5231(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2F00B),
				.b1(W2F01B),
				.b2(W2F02B),
				.b3(W2F10B),
				.b4(W2F11B),
				.b5(W2F12B),
				.b6(W2F20B),
				.b7(W2F21B),
				.b8(W2F22B),
				.c(c2B20F)
);

ninexnine_unit ninexnine_unit_5232(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2F00C),
				.b1(W2F01C),
				.b2(W2F02C),
				.b3(W2F10C),
				.b4(W2F11C),
				.b5(W2F12C),
				.b6(W2F20C),
				.b7(W2F21C),
				.b8(W2F22C),
				.c(c2C20F)
);

ninexnine_unit ninexnine_unit_5233(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2F00D),
				.b1(W2F01D),
				.b2(W2F02D),
				.b3(W2F10D),
				.b4(W2F11D),
				.b5(W2F12D),
				.b6(W2F20D),
				.b7(W2F21D),
				.b8(W2F22D),
				.c(c2D20F)
);

ninexnine_unit ninexnine_unit_5234(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2F00E),
				.b1(W2F01E),
				.b2(W2F02E),
				.b3(W2F10E),
				.b4(W2F11E),
				.b5(W2F12E),
				.b6(W2F20E),
				.b7(W2F21E),
				.b8(W2F22E),
				.c(c2E20F)
);

ninexnine_unit ninexnine_unit_5235(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2F00F),
				.b1(W2F01F),
				.b2(W2F02F),
				.b3(W2F10F),
				.b4(W2F11F),
				.b5(W2F12F),
				.b6(W2F20F),
				.b7(W2F21F),
				.b8(W2F22F),
				.c(c2F20F)
);

assign C220F=c2020F+c2120F+c2220F+c2320F+c2420F+c2520F+c2620F+c2720F+c2820F+c2920F+c2A20F+c2B20F+c2C20F+c2D20F+c2E20F+c2F20F;
assign A220F=(C220F>=0)?1:0;

assign P320F=A220F;

ninexnine_unit ninexnine_unit_5236(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2021F)
);

ninexnine_unit ninexnine_unit_5237(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2121F)
);

ninexnine_unit ninexnine_unit_5238(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2221F)
);

ninexnine_unit ninexnine_unit_5239(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2321F)
);

ninexnine_unit ninexnine_unit_5240(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2421F)
);

ninexnine_unit ninexnine_unit_5241(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2521F)
);

ninexnine_unit ninexnine_unit_5242(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2621F)
);

ninexnine_unit ninexnine_unit_5243(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2721F)
);

ninexnine_unit ninexnine_unit_5244(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2F008),
				.b1(W2F018),
				.b2(W2F028),
				.b3(W2F108),
				.b4(W2F118),
				.b5(W2F128),
				.b6(W2F208),
				.b7(W2F218),
				.b8(W2F228),
				.c(c2821F)
);

ninexnine_unit ninexnine_unit_5245(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2F009),
				.b1(W2F019),
				.b2(W2F029),
				.b3(W2F109),
				.b4(W2F119),
				.b5(W2F129),
				.b6(W2F209),
				.b7(W2F219),
				.b8(W2F229),
				.c(c2921F)
);

ninexnine_unit ninexnine_unit_5246(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2F00A),
				.b1(W2F01A),
				.b2(W2F02A),
				.b3(W2F10A),
				.b4(W2F11A),
				.b5(W2F12A),
				.b6(W2F20A),
				.b7(W2F21A),
				.b8(W2F22A),
				.c(c2A21F)
);

ninexnine_unit ninexnine_unit_5247(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2F00B),
				.b1(W2F01B),
				.b2(W2F02B),
				.b3(W2F10B),
				.b4(W2F11B),
				.b5(W2F12B),
				.b6(W2F20B),
				.b7(W2F21B),
				.b8(W2F22B),
				.c(c2B21F)
);

ninexnine_unit ninexnine_unit_5248(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2F00C),
				.b1(W2F01C),
				.b2(W2F02C),
				.b3(W2F10C),
				.b4(W2F11C),
				.b5(W2F12C),
				.b6(W2F20C),
				.b7(W2F21C),
				.b8(W2F22C),
				.c(c2C21F)
);

ninexnine_unit ninexnine_unit_5249(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2F00D),
				.b1(W2F01D),
				.b2(W2F02D),
				.b3(W2F10D),
				.b4(W2F11D),
				.b5(W2F12D),
				.b6(W2F20D),
				.b7(W2F21D),
				.b8(W2F22D),
				.c(c2D21F)
);

ninexnine_unit ninexnine_unit_5250(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2F00E),
				.b1(W2F01E),
				.b2(W2F02E),
				.b3(W2F10E),
				.b4(W2F11E),
				.b5(W2F12E),
				.b6(W2F20E),
				.b7(W2F21E),
				.b8(W2F22E),
				.c(c2E21F)
);

ninexnine_unit ninexnine_unit_5251(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2F00F),
				.b1(W2F01F),
				.b2(W2F02F),
				.b3(W2F10F),
				.b4(W2F11F),
				.b5(W2F12F),
				.b6(W2F20F),
				.b7(W2F21F),
				.b8(W2F22F),
				.c(c2F21F)
);

assign C221F=c2021F+c2121F+c2221F+c2321F+c2421F+c2521F+c2621F+c2721F+c2821F+c2921F+c2A21F+c2B21F+c2C21F+c2D21F+c2E21F+c2F21F;
assign A221F=(C221F>=0)?1:0;

assign P321F=A221F;

ninexnine_unit ninexnine_unit_5252(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2F000),
				.b1(W2F010),
				.b2(W2F020),
				.b3(W2F100),
				.b4(W2F110),
				.b5(W2F120),
				.b6(W2F200),
				.b7(W2F210),
				.b8(W2F220),
				.c(c2022F)
);

ninexnine_unit ninexnine_unit_5253(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2F001),
				.b1(W2F011),
				.b2(W2F021),
				.b3(W2F101),
				.b4(W2F111),
				.b5(W2F121),
				.b6(W2F201),
				.b7(W2F211),
				.b8(W2F221),
				.c(c2122F)
);

ninexnine_unit ninexnine_unit_5254(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2F002),
				.b1(W2F012),
				.b2(W2F022),
				.b3(W2F102),
				.b4(W2F112),
				.b5(W2F122),
				.b6(W2F202),
				.b7(W2F212),
				.b8(W2F222),
				.c(c2222F)
);

ninexnine_unit ninexnine_unit_5255(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2F003),
				.b1(W2F013),
				.b2(W2F023),
				.b3(W2F103),
				.b4(W2F113),
				.b5(W2F123),
				.b6(W2F203),
				.b7(W2F213),
				.b8(W2F223),
				.c(c2322F)
);

ninexnine_unit ninexnine_unit_5256(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2F004),
				.b1(W2F014),
				.b2(W2F024),
				.b3(W2F104),
				.b4(W2F114),
				.b5(W2F124),
				.b6(W2F204),
				.b7(W2F214),
				.b8(W2F224),
				.c(c2422F)
);

ninexnine_unit ninexnine_unit_5257(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2F005),
				.b1(W2F015),
				.b2(W2F025),
				.b3(W2F105),
				.b4(W2F115),
				.b5(W2F125),
				.b6(W2F205),
				.b7(W2F215),
				.b8(W2F225),
				.c(c2522F)
);

ninexnine_unit ninexnine_unit_5258(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2F006),
				.b1(W2F016),
				.b2(W2F026),
				.b3(W2F106),
				.b4(W2F116),
				.b5(W2F126),
				.b6(W2F206),
				.b7(W2F216),
				.b8(W2F226),
				.c(c2622F)
);

ninexnine_unit ninexnine_unit_5259(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2F007),
				.b1(W2F017),
				.b2(W2F027),
				.b3(W2F107),
				.b4(W2F117),
				.b5(W2F127),
				.b6(W2F207),
				.b7(W2F217),
				.b8(W2F227),
				.c(c2722F)
);

ninexnine_unit ninexnine_unit_5260(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2F008),
				.b1(W2F018),
				.b2(W2F028),
				.b3(W2F108),
				.b4(W2F118),
				.b5(W2F128),
				.b6(W2F208),
				.b7(W2F218),
				.b8(W2F228),
				.c(c2822F)
);

ninexnine_unit ninexnine_unit_5261(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2F009),
				.b1(W2F019),
				.b2(W2F029),
				.b3(W2F109),
				.b4(W2F119),
				.b5(W2F129),
				.b6(W2F209),
				.b7(W2F219),
				.b8(W2F229),
				.c(c2922F)
);

ninexnine_unit ninexnine_unit_5262(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2F00A),
				.b1(W2F01A),
				.b2(W2F02A),
				.b3(W2F10A),
				.b4(W2F11A),
				.b5(W2F12A),
				.b6(W2F20A),
				.b7(W2F21A),
				.b8(W2F22A),
				.c(c2A22F)
);

ninexnine_unit ninexnine_unit_5263(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2F00B),
				.b1(W2F01B),
				.b2(W2F02B),
				.b3(W2F10B),
				.b4(W2F11B),
				.b5(W2F12B),
				.b6(W2F20B),
				.b7(W2F21B),
				.b8(W2F22B),
				.c(c2B22F)
);

ninexnine_unit ninexnine_unit_5264(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2F00C),
				.b1(W2F01C),
				.b2(W2F02C),
				.b3(W2F10C),
				.b4(W2F11C),
				.b5(W2F12C),
				.b6(W2F20C),
				.b7(W2F21C),
				.b8(W2F22C),
				.c(c2C22F)
);

ninexnine_unit ninexnine_unit_5265(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2F00D),
				.b1(W2F01D),
				.b2(W2F02D),
				.b3(W2F10D),
				.b4(W2F11D),
				.b5(W2F12D),
				.b6(W2F20D),
				.b7(W2F21D),
				.b8(W2F22D),
				.c(c2D22F)
);

ninexnine_unit ninexnine_unit_5266(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2F00E),
				.b1(W2F01E),
				.b2(W2F02E),
				.b3(W2F10E),
				.b4(W2F11E),
				.b5(W2F12E),
				.b6(W2F20E),
				.b7(W2F21E),
				.b8(W2F22E),
				.c(c2E22F)
);

ninexnine_unit ninexnine_unit_5267(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2F00F),
				.b1(W2F01F),
				.b2(W2F02F),
				.b3(W2F10F),
				.b4(W2F11F),
				.b5(W2F12F),
				.b6(W2F20F),
				.b7(W2F21F),
				.b8(W2F22F),
				.c(c2F22F)
);

assign C222F=c2022F+c2122F+c2222F+c2322F+c2422F+c2522F+c2622F+c2722F+c2822F+c2922F+c2A22F+c2B22F+c2C22F+c2D22F+c2E22F+c2F22F;
assign A222F=(C222F>=0)?1:0;

assign P322F=A222F;

ninexnine_unit ninexnine_unit_5268(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2G000),
				.b1(W2G010),
				.b2(W2G020),
				.b3(W2G100),
				.b4(W2G110),
				.b5(W2G120),
				.b6(W2G200),
				.b7(W2G210),
				.b8(W2G220),
				.c(c2000G)
);

ninexnine_unit ninexnine_unit_5269(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2G001),
				.b1(W2G011),
				.b2(W2G021),
				.b3(W2G101),
				.b4(W2G111),
				.b5(W2G121),
				.b6(W2G201),
				.b7(W2G211),
				.b8(W2G221),
				.c(c2100G)
);

ninexnine_unit ninexnine_unit_5270(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2G002),
				.b1(W2G012),
				.b2(W2G022),
				.b3(W2G102),
				.b4(W2G112),
				.b5(W2G122),
				.b6(W2G202),
				.b7(W2G212),
				.b8(W2G222),
				.c(c2200G)
);

ninexnine_unit ninexnine_unit_5271(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2G003),
				.b1(W2G013),
				.b2(W2G023),
				.b3(W2G103),
				.b4(W2G113),
				.b5(W2G123),
				.b6(W2G203),
				.b7(W2G213),
				.b8(W2G223),
				.c(c2300G)
);

ninexnine_unit ninexnine_unit_5272(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2G004),
				.b1(W2G014),
				.b2(W2G024),
				.b3(W2G104),
				.b4(W2G114),
				.b5(W2G124),
				.b6(W2G204),
				.b7(W2G214),
				.b8(W2G224),
				.c(c2400G)
);

ninexnine_unit ninexnine_unit_5273(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2G005),
				.b1(W2G015),
				.b2(W2G025),
				.b3(W2G105),
				.b4(W2G115),
				.b5(W2G125),
				.b6(W2G205),
				.b7(W2G215),
				.b8(W2G225),
				.c(c2500G)
);

ninexnine_unit ninexnine_unit_5274(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2G006),
				.b1(W2G016),
				.b2(W2G026),
				.b3(W2G106),
				.b4(W2G116),
				.b5(W2G126),
				.b6(W2G206),
				.b7(W2G216),
				.b8(W2G226),
				.c(c2600G)
);

ninexnine_unit ninexnine_unit_5275(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2G007),
				.b1(W2G017),
				.b2(W2G027),
				.b3(W2G107),
				.b4(W2G117),
				.b5(W2G127),
				.b6(W2G207),
				.b7(W2G217),
				.b8(W2G227),
				.c(c2700G)
);

ninexnine_unit ninexnine_unit_5276(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2G008),
				.b1(W2G018),
				.b2(W2G028),
				.b3(W2G108),
				.b4(W2G118),
				.b5(W2G128),
				.b6(W2G208),
				.b7(W2G218),
				.b8(W2G228),
				.c(c2800G)
);

ninexnine_unit ninexnine_unit_5277(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2G009),
				.b1(W2G019),
				.b2(W2G029),
				.b3(W2G109),
				.b4(W2G119),
				.b5(W2G129),
				.b6(W2G209),
				.b7(W2G219),
				.b8(W2G229),
				.c(c2900G)
);

ninexnine_unit ninexnine_unit_5278(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2G00A),
				.b1(W2G01A),
				.b2(W2G02A),
				.b3(W2G10A),
				.b4(W2G11A),
				.b5(W2G12A),
				.b6(W2G20A),
				.b7(W2G21A),
				.b8(W2G22A),
				.c(c2A00G)
);

ninexnine_unit ninexnine_unit_5279(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2G00B),
				.b1(W2G01B),
				.b2(W2G02B),
				.b3(W2G10B),
				.b4(W2G11B),
				.b5(W2G12B),
				.b6(W2G20B),
				.b7(W2G21B),
				.b8(W2G22B),
				.c(c2B00G)
);

ninexnine_unit ninexnine_unit_5280(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2G00C),
				.b1(W2G01C),
				.b2(W2G02C),
				.b3(W2G10C),
				.b4(W2G11C),
				.b5(W2G12C),
				.b6(W2G20C),
				.b7(W2G21C),
				.b8(W2G22C),
				.c(c2C00G)
);

ninexnine_unit ninexnine_unit_5281(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2G00D),
				.b1(W2G01D),
				.b2(W2G02D),
				.b3(W2G10D),
				.b4(W2G11D),
				.b5(W2G12D),
				.b6(W2G20D),
				.b7(W2G21D),
				.b8(W2G22D),
				.c(c2D00G)
);

ninexnine_unit ninexnine_unit_5282(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2G00E),
				.b1(W2G01E),
				.b2(W2G02E),
				.b3(W2G10E),
				.b4(W2G11E),
				.b5(W2G12E),
				.b6(W2G20E),
				.b7(W2G21E),
				.b8(W2G22E),
				.c(c2E00G)
);

ninexnine_unit ninexnine_unit_5283(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2G00F),
				.b1(W2G01F),
				.b2(W2G02F),
				.b3(W2G10F),
				.b4(W2G11F),
				.b5(W2G12F),
				.b6(W2G20F),
				.b7(W2G21F),
				.b8(W2G22F),
				.c(c2F00G)
);

assign C200G=c2000G+c2100G+c2200G+c2300G+c2400G+c2500G+c2600G+c2700G+c2800G+c2900G+c2A00G+c2B00G+c2C00G+c2D00G+c2E00G+c2F00G;
assign A200G=(C200G>=0)?1:0;

assign P300G=A200G;

ninexnine_unit ninexnine_unit_5284(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2G000),
				.b1(W2G010),
				.b2(W2G020),
				.b3(W2G100),
				.b4(W2G110),
				.b5(W2G120),
				.b6(W2G200),
				.b7(W2G210),
				.b8(W2G220),
				.c(c2001G)
);

ninexnine_unit ninexnine_unit_5285(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2G001),
				.b1(W2G011),
				.b2(W2G021),
				.b3(W2G101),
				.b4(W2G111),
				.b5(W2G121),
				.b6(W2G201),
				.b7(W2G211),
				.b8(W2G221),
				.c(c2101G)
);

ninexnine_unit ninexnine_unit_5286(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2G002),
				.b1(W2G012),
				.b2(W2G022),
				.b3(W2G102),
				.b4(W2G112),
				.b5(W2G122),
				.b6(W2G202),
				.b7(W2G212),
				.b8(W2G222),
				.c(c2201G)
);

ninexnine_unit ninexnine_unit_5287(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2G003),
				.b1(W2G013),
				.b2(W2G023),
				.b3(W2G103),
				.b4(W2G113),
				.b5(W2G123),
				.b6(W2G203),
				.b7(W2G213),
				.b8(W2G223),
				.c(c2301G)
);

ninexnine_unit ninexnine_unit_5288(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2G004),
				.b1(W2G014),
				.b2(W2G024),
				.b3(W2G104),
				.b4(W2G114),
				.b5(W2G124),
				.b6(W2G204),
				.b7(W2G214),
				.b8(W2G224),
				.c(c2401G)
);

ninexnine_unit ninexnine_unit_5289(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2G005),
				.b1(W2G015),
				.b2(W2G025),
				.b3(W2G105),
				.b4(W2G115),
				.b5(W2G125),
				.b6(W2G205),
				.b7(W2G215),
				.b8(W2G225),
				.c(c2501G)
);

ninexnine_unit ninexnine_unit_5290(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2G006),
				.b1(W2G016),
				.b2(W2G026),
				.b3(W2G106),
				.b4(W2G116),
				.b5(W2G126),
				.b6(W2G206),
				.b7(W2G216),
				.b8(W2G226),
				.c(c2601G)
);

ninexnine_unit ninexnine_unit_5291(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2G007),
				.b1(W2G017),
				.b2(W2G027),
				.b3(W2G107),
				.b4(W2G117),
				.b5(W2G127),
				.b6(W2G207),
				.b7(W2G217),
				.b8(W2G227),
				.c(c2701G)
);

ninexnine_unit ninexnine_unit_5292(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2G008),
				.b1(W2G018),
				.b2(W2G028),
				.b3(W2G108),
				.b4(W2G118),
				.b5(W2G128),
				.b6(W2G208),
				.b7(W2G218),
				.b8(W2G228),
				.c(c2801G)
);

ninexnine_unit ninexnine_unit_5293(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2G009),
				.b1(W2G019),
				.b2(W2G029),
				.b3(W2G109),
				.b4(W2G119),
				.b5(W2G129),
				.b6(W2G209),
				.b7(W2G219),
				.b8(W2G229),
				.c(c2901G)
);

ninexnine_unit ninexnine_unit_5294(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2G00A),
				.b1(W2G01A),
				.b2(W2G02A),
				.b3(W2G10A),
				.b4(W2G11A),
				.b5(W2G12A),
				.b6(W2G20A),
				.b7(W2G21A),
				.b8(W2G22A),
				.c(c2A01G)
);

ninexnine_unit ninexnine_unit_5295(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2G00B),
				.b1(W2G01B),
				.b2(W2G02B),
				.b3(W2G10B),
				.b4(W2G11B),
				.b5(W2G12B),
				.b6(W2G20B),
				.b7(W2G21B),
				.b8(W2G22B),
				.c(c2B01G)
);

ninexnine_unit ninexnine_unit_5296(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2G00C),
				.b1(W2G01C),
				.b2(W2G02C),
				.b3(W2G10C),
				.b4(W2G11C),
				.b5(W2G12C),
				.b6(W2G20C),
				.b7(W2G21C),
				.b8(W2G22C),
				.c(c2C01G)
);

ninexnine_unit ninexnine_unit_5297(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2G00D),
				.b1(W2G01D),
				.b2(W2G02D),
				.b3(W2G10D),
				.b4(W2G11D),
				.b5(W2G12D),
				.b6(W2G20D),
				.b7(W2G21D),
				.b8(W2G22D),
				.c(c2D01G)
);

ninexnine_unit ninexnine_unit_5298(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2G00E),
				.b1(W2G01E),
				.b2(W2G02E),
				.b3(W2G10E),
				.b4(W2G11E),
				.b5(W2G12E),
				.b6(W2G20E),
				.b7(W2G21E),
				.b8(W2G22E),
				.c(c2E01G)
);

ninexnine_unit ninexnine_unit_5299(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2G00F),
				.b1(W2G01F),
				.b2(W2G02F),
				.b3(W2G10F),
				.b4(W2G11F),
				.b5(W2G12F),
				.b6(W2G20F),
				.b7(W2G21F),
				.b8(W2G22F),
				.c(c2F01G)
);

assign C201G=c2001G+c2101G+c2201G+c2301G+c2401G+c2501G+c2601G+c2701G+c2801G+c2901G+c2A01G+c2B01G+c2C01G+c2D01G+c2E01G+c2F01G;
assign A201G=(C201G>=0)?1:0;

assign P301G=A201G;

ninexnine_unit ninexnine_unit_5300(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2G000),
				.b1(W2G010),
				.b2(W2G020),
				.b3(W2G100),
				.b4(W2G110),
				.b5(W2G120),
				.b6(W2G200),
				.b7(W2G210),
				.b8(W2G220),
				.c(c2002G)
);

ninexnine_unit ninexnine_unit_5301(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2G001),
				.b1(W2G011),
				.b2(W2G021),
				.b3(W2G101),
				.b4(W2G111),
				.b5(W2G121),
				.b6(W2G201),
				.b7(W2G211),
				.b8(W2G221),
				.c(c2102G)
);

ninexnine_unit ninexnine_unit_5302(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2G002),
				.b1(W2G012),
				.b2(W2G022),
				.b3(W2G102),
				.b4(W2G112),
				.b5(W2G122),
				.b6(W2G202),
				.b7(W2G212),
				.b8(W2G222),
				.c(c2202G)
);

ninexnine_unit ninexnine_unit_5303(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2G003),
				.b1(W2G013),
				.b2(W2G023),
				.b3(W2G103),
				.b4(W2G113),
				.b5(W2G123),
				.b6(W2G203),
				.b7(W2G213),
				.b8(W2G223),
				.c(c2302G)
);

ninexnine_unit ninexnine_unit_5304(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2G004),
				.b1(W2G014),
				.b2(W2G024),
				.b3(W2G104),
				.b4(W2G114),
				.b5(W2G124),
				.b6(W2G204),
				.b7(W2G214),
				.b8(W2G224),
				.c(c2402G)
);

ninexnine_unit ninexnine_unit_5305(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2G005),
				.b1(W2G015),
				.b2(W2G025),
				.b3(W2G105),
				.b4(W2G115),
				.b5(W2G125),
				.b6(W2G205),
				.b7(W2G215),
				.b8(W2G225),
				.c(c2502G)
);

ninexnine_unit ninexnine_unit_5306(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2G006),
				.b1(W2G016),
				.b2(W2G026),
				.b3(W2G106),
				.b4(W2G116),
				.b5(W2G126),
				.b6(W2G206),
				.b7(W2G216),
				.b8(W2G226),
				.c(c2602G)
);

ninexnine_unit ninexnine_unit_5307(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2G007),
				.b1(W2G017),
				.b2(W2G027),
				.b3(W2G107),
				.b4(W2G117),
				.b5(W2G127),
				.b6(W2G207),
				.b7(W2G217),
				.b8(W2G227),
				.c(c2702G)
);

ninexnine_unit ninexnine_unit_5308(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2G008),
				.b1(W2G018),
				.b2(W2G028),
				.b3(W2G108),
				.b4(W2G118),
				.b5(W2G128),
				.b6(W2G208),
				.b7(W2G218),
				.b8(W2G228),
				.c(c2802G)
);

ninexnine_unit ninexnine_unit_5309(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2G009),
				.b1(W2G019),
				.b2(W2G029),
				.b3(W2G109),
				.b4(W2G119),
				.b5(W2G129),
				.b6(W2G209),
				.b7(W2G219),
				.b8(W2G229),
				.c(c2902G)
);

ninexnine_unit ninexnine_unit_5310(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2G00A),
				.b1(W2G01A),
				.b2(W2G02A),
				.b3(W2G10A),
				.b4(W2G11A),
				.b5(W2G12A),
				.b6(W2G20A),
				.b7(W2G21A),
				.b8(W2G22A),
				.c(c2A02G)
);

ninexnine_unit ninexnine_unit_5311(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2G00B),
				.b1(W2G01B),
				.b2(W2G02B),
				.b3(W2G10B),
				.b4(W2G11B),
				.b5(W2G12B),
				.b6(W2G20B),
				.b7(W2G21B),
				.b8(W2G22B),
				.c(c2B02G)
);

ninexnine_unit ninexnine_unit_5312(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2G00C),
				.b1(W2G01C),
				.b2(W2G02C),
				.b3(W2G10C),
				.b4(W2G11C),
				.b5(W2G12C),
				.b6(W2G20C),
				.b7(W2G21C),
				.b8(W2G22C),
				.c(c2C02G)
);

ninexnine_unit ninexnine_unit_5313(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2G00D),
				.b1(W2G01D),
				.b2(W2G02D),
				.b3(W2G10D),
				.b4(W2G11D),
				.b5(W2G12D),
				.b6(W2G20D),
				.b7(W2G21D),
				.b8(W2G22D),
				.c(c2D02G)
);

ninexnine_unit ninexnine_unit_5314(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2G00E),
				.b1(W2G01E),
				.b2(W2G02E),
				.b3(W2G10E),
				.b4(W2G11E),
				.b5(W2G12E),
				.b6(W2G20E),
				.b7(W2G21E),
				.b8(W2G22E),
				.c(c2E02G)
);

ninexnine_unit ninexnine_unit_5315(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2G00F),
				.b1(W2G01F),
				.b2(W2G02F),
				.b3(W2G10F),
				.b4(W2G11F),
				.b5(W2G12F),
				.b6(W2G20F),
				.b7(W2G21F),
				.b8(W2G22F),
				.c(c2F02G)
);

assign C202G=c2002G+c2102G+c2202G+c2302G+c2402G+c2502G+c2602G+c2702G+c2802G+c2902G+c2A02G+c2B02G+c2C02G+c2D02G+c2E02G+c2F02G;
assign A202G=(C202G>=0)?1:0;

assign P302G=A202G;

ninexnine_unit ninexnine_unit_5316(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2G000),
				.b1(W2G010),
				.b2(W2G020),
				.b3(W2G100),
				.b4(W2G110),
				.b5(W2G120),
				.b6(W2G200),
				.b7(W2G210),
				.b8(W2G220),
				.c(c2010G)
);

ninexnine_unit ninexnine_unit_5317(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2G001),
				.b1(W2G011),
				.b2(W2G021),
				.b3(W2G101),
				.b4(W2G111),
				.b5(W2G121),
				.b6(W2G201),
				.b7(W2G211),
				.b8(W2G221),
				.c(c2110G)
);

ninexnine_unit ninexnine_unit_5318(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2G002),
				.b1(W2G012),
				.b2(W2G022),
				.b3(W2G102),
				.b4(W2G112),
				.b5(W2G122),
				.b6(W2G202),
				.b7(W2G212),
				.b8(W2G222),
				.c(c2210G)
);

ninexnine_unit ninexnine_unit_5319(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2G003),
				.b1(W2G013),
				.b2(W2G023),
				.b3(W2G103),
				.b4(W2G113),
				.b5(W2G123),
				.b6(W2G203),
				.b7(W2G213),
				.b8(W2G223),
				.c(c2310G)
);

ninexnine_unit ninexnine_unit_5320(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2G004),
				.b1(W2G014),
				.b2(W2G024),
				.b3(W2G104),
				.b4(W2G114),
				.b5(W2G124),
				.b6(W2G204),
				.b7(W2G214),
				.b8(W2G224),
				.c(c2410G)
);

ninexnine_unit ninexnine_unit_5321(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2G005),
				.b1(W2G015),
				.b2(W2G025),
				.b3(W2G105),
				.b4(W2G115),
				.b5(W2G125),
				.b6(W2G205),
				.b7(W2G215),
				.b8(W2G225),
				.c(c2510G)
);

ninexnine_unit ninexnine_unit_5322(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2G006),
				.b1(W2G016),
				.b2(W2G026),
				.b3(W2G106),
				.b4(W2G116),
				.b5(W2G126),
				.b6(W2G206),
				.b7(W2G216),
				.b8(W2G226),
				.c(c2610G)
);

ninexnine_unit ninexnine_unit_5323(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2G007),
				.b1(W2G017),
				.b2(W2G027),
				.b3(W2G107),
				.b4(W2G117),
				.b5(W2G127),
				.b6(W2G207),
				.b7(W2G217),
				.b8(W2G227),
				.c(c2710G)
);

ninexnine_unit ninexnine_unit_5324(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2G008),
				.b1(W2G018),
				.b2(W2G028),
				.b3(W2G108),
				.b4(W2G118),
				.b5(W2G128),
				.b6(W2G208),
				.b7(W2G218),
				.b8(W2G228),
				.c(c2810G)
);

ninexnine_unit ninexnine_unit_5325(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2G009),
				.b1(W2G019),
				.b2(W2G029),
				.b3(W2G109),
				.b4(W2G119),
				.b5(W2G129),
				.b6(W2G209),
				.b7(W2G219),
				.b8(W2G229),
				.c(c2910G)
);

ninexnine_unit ninexnine_unit_5326(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2G00A),
				.b1(W2G01A),
				.b2(W2G02A),
				.b3(W2G10A),
				.b4(W2G11A),
				.b5(W2G12A),
				.b6(W2G20A),
				.b7(W2G21A),
				.b8(W2G22A),
				.c(c2A10G)
);

ninexnine_unit ninexnine_unit_5327(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2G00B),
				.b1(W2G01B),
				.b2(W2G02B),
				.b3(W2G10B),
				.b4(W2G11B),
				.b5(W2G12B),
				.b6(W2G20B),
				.b7(W2G21B),
				.b8(W2G22B),
				.c(c2B10G)
);

ninexnine_unit ninexnine_unit_5328(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2G00C),
				.b1(W2G01C),
				.b2(W2G02C),
				.b3(W2G10C),
				.b4(W2G11C),
				.b5(W2G12C),
				.b6(W2G20C),
				.b7(W2G21C),
				.b8(W2G22C),
				.c(c2C10G)
);

ninexnine_unit ninexnine_unit_5329(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2G00D),
				.b1(W2G01D),
				.b2(W2G02D),
				.b3(W2G10D),
				.b4(W2G11D),
				.b5(W2G12D),
				.b6(W2G20D),
				.b7(W2G21D),
				.b8(W2G22D),
				.c(c2D10G)
);

ninexnine_unit ninexnine_unit_5330(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2G00E),
				.b1(W2G01E),
				.b2(W2G02E),
				.b3(W2G10E),
				.b4(W2G11E),
				.b5(W2G12E),
				.b6(W2G20E),
				.b7(W2G21E),
				.b8(W2G22E),
				.c(c2E10G)
);

ninexnine_unit ninexnine_unit_5331(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2G00F),
				.b1(W2G01F),
				.b2(W2G02F),
				.b3(W2G10F),
				.b4(W2G11F),
				.b5(W2G12F),
				.b6(W2G20F),
				.b7(W2G21F),
				.b8(W2G22F),
				.c(c2F10G)
);

assign C210G=c2010G+c2110G+c2210G+c2310G+c2410G+c2510G+c2610G+c2710G+c2810G+c2910G+c2A10G+c2B10G+c2C10G+c2D10G+c2E10G+c2F10G;
assign A210G=(C210G>=0)?1:0;

assign P310G=A210G;

ninexnine_unit ninexnine_unit_5332(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2G000),
				.b1(W2G010),
				.b2(W2G020),
				.b3(W2G100),
				.b4(W2G110),
				.b5(W2G120),
				.b6(W2G200),
				.b7(W2G210),
				.b8(W2G220),
				.c(c2011G)
);

ninexnine_unit ninexnine_unit_5333(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2G001),
				.b1(W2G011),
				.b2(W2G021),
				.b3(W2G101),
				.b4(W2G111),
				.b5(W2G121),
				.b6(W2G201),
				.b7(W2G211),
				.b8(W2G221),
				.c(c2111G)
);

ninexnine_unit ninexnine_unit_5334(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2G002),
				.b1(W2G012),
				.b2(W2G022),
				.b3(W2G102),
				.b4(W2G112),
				.b5(W2G122),
				.b6(W2G202),
				.b7(W2G212),
				.b8(W2G222),
				.c(c2211G)
);

ninexnine_unit ninexnine_unit_5335(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2G003),
				.b1(W2G013),
				.b2(W2G023),
				.b3(W2G103),
				.b4(W2G113),
				.b5(W2G123),
				.b6(W2G203),
				.b7(W2G213),
				.b8(W2G223),
				.c(c2311G)
);

ninexnine_unit ninexnine_unit_5336(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2G004),
				.b1(W2G014),
				.b2(W2G024),
				.b3(W2G104),
				.b4(W2G114),
				.b5(W2G124),
				.b6(W2G204),
				.b7(W2G214),
				.b8(W2G224),
				.c(c2411G)
);

ninexnine_unit ninexnine_unit_5337(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2G005),
				.b1(W2G015),
				.b2(W2G025),
				.b3(W2G105),
				.b4(W2G115),
				.b5(W2G125),
				.b6(W2G205),
				.b7(W2G215),
				.b8(W2G225),
				.c(c2511G)
);

ninexnine_unit ninexnine_unit_5338(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2G006),
				.b1(W2G016),
				.b2(W2G026),
				.b3(W2G106),
				.b4(W2G116),
				.b5(W2G126),
				.b6(W2G206),
				.b7(W2G216),
				.b8(W2G226),
				.c(c2611G)
);

ninexnine_unit ninexnine_unit_5339(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2G007),
				.b1(W2G017),
				.b2(W2G027),
				.b3(W2G107),
				.b4(W2G117),
				.b5(W2G127),
				.b6(W2G207),
				.b7(W2G217),
				.b8(W2G227),
				.c(c2711G)
);

ninexnine_unit ninexnine_unit_5340(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2G008),
				.b1(W2G018),
				.b2(W2G028),
				.b3(W2G108),
				.b4(W2G118),
				.b5(W2G128),
				.b6(W2G208),
				.b7(W2G218),
				.b8(W2G228),
				.c(c2811G)
);

ninexnine_unit ninexnine_unit_5341(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2G009),
				.b1(W2G019),
				.b2(W2G029),
				.b3(W2G109),
				.b4(W2G119),
				.b5(W2G129),
				.b6(W2G209),
				.b7(W2G219),
				.b8(W2G229),
				.c(c2911G)
);

ninexnine_unit ninexnine_unit_5342(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2G00A),
				.b1(W2G01A),
				.b2(W2G02A),
				.b3(W2G10A),
				.b4(W2G11A),
				.b5(W2G12A),
				.b6(W2G20A),
				.b7(W2G21A),
				.b8(W2G22A),
				.c(c2A11G)
);

ninexnine_unit ninexnine_unit_5343(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2G00B),
				.b1(W2G01B),
				.b2(W2G02B),
				.b3(W2G10B),
				.b4(W2G11B),
				.b5(W2G12B),
				.b6(W2G20B),
				.b7(W2G21B),
				.b8(W2G22B),
				.c(c2B11G)
);

ninexnine_unit ninexnine_unit_5344(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2G00C),
				.b1(W2G01C),
				.b2(W2G02C),
				.b3(W2G10C),
				.b4(W2G11C),
				.b5(W2G12C),
				.b6(W2G20C),
				.b7(W2G21C),
				.b8(W2G22C),
				.c(c2C11G)
);

ninexnine_unit ninexnine_unit_5345(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2G00D),
				.b1(W2G01D),
				.b2(W2G02D),
				.b3(W2G10D),
				.b4(W2G11D),
				.b5(W2G12D),
				.b6(W2G20D),
				.b7(W2G21D),
				.b8(W2G22D),
				.c(c2D11G)
);

ninexnine_unit ninexnine_unit_5346(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2G00E),
				.b1(W2G01E),
				.b2(W2G02E),
				.b3(W2G10E),
				.b4(W2G11E),
				.b5(W2G12E),
				.b6(W2G20E),
				.b7(W2G21E),
				.b8(W2G22E),
				.c(c2E11G)
);

ninexnine_unit ninexnine_unit_5347(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2G00F),
				.b1(W2G01F),
				.b2(W2G02F),
				.b3(W2G10F),
				.b4(W2G11F),
				.b5(W2G12F),
				.b6(W2G20F),
				.b7(W2G21F),
				.b8(W2G22F),
				.c(c2F11G)
);

assign C211G=c2011G+c2111G+c2211G+c2311G+c2411G+c2511G+c2611G+c2711G+c2811G+c2911G+c2A11G+c2B11G+c2C11G+c2D11G+c2E11G+c2F11G;
assign A211G=(C211G>=0)?1:0;

assign P311G=A211G;

ninexnine_unit ninexnine_unit_5348(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2G000),
				.b1(W2G010),
				.b2(W2G020),
				.b3(W2G100),
				.b4(W2G110),
				.b5(W2G120),
				.b6(W2G200),
				.b7(W2G210),
				.b8(W2G220),
				.c(c2012G)
);

ninexnine_unit ninexnine_unit_5349(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2G001),
				.b1(W2G011),
				.b2(W2G021),
				.b3(W2G101),
				.b4(W2G111),
				.b5(W2G121),
				.b6(W2G201),
				.b7(W2G211),
				.b8(W2G221),
				.c(c2112G)
);

ninexnine_unit ninexnine_unit_5350(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2G002),
				.b1(W2G012),
				.b2(W2G022),
				.b3(W2G102),
				.b4(W2G112),
				.b5(W2G122),
				.b6(W2G202),
				.b7(W2G212),
				.b8(W2G222),
				.c(c2212G)
);

ninexnine_unit ninexnine_unit_5351(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2G003),
				.b1(W2G013),
				.b2(W2G023),
				.b3(W2G103),
				.b4(W2G113),
				.b5(W2G123),
				.b6(W2G203),
				.b7(W2G213),
				.b8(W2G223),
				.c(c2312G)
);

ninexnine_unit ninexnine_unit_5352(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2G004),
				.b1(W2G014),
				.b2(W2G024),
				.b3(W2G104),
				.b4(W2G114),
				.b5(W2G124),
				.b6(W2G204),
				.b7(W2G214),
				.b8(W2G224),
				.c(c2412G)
);

ninexnine_unit ninexnine_unit_5353(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2G005),
				.b1(W2G015),
				.b2(W2G025),
				.b3(W2G105),
				.b4(W2G115),
				.b5(W2G125),
				.b6(W2G205),
				.b7(W2G215),
				.b8(W2G225),
				.c(c2512G)
);

ninexnine_unit ninexnine_unit_5354(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2G006),
				.b1(W2G016),
				.b2(W2G026),
				.b3(W2G106),
				.b4(W2G116),
				.b5(W2G126),
				.b6(W2G206),
				.b7(W2G216),
				.b8(W2G226),
				.c(c2612G)
);

ninexnine_unit ninexnine_unit_5355(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2G007),
				.b1(W2G017),
				.b2(W2G027),
				.b3(W2G107),
				.b4(W2G117),
				.b5(W2G127),
				.b6(W2G207),
				.b7(W2G217),
				.b8(W2G227),
				.c(c2712G)
);

ninexnine_unit ninexnine_unit_5356(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2G008),
				.b1(W2G018),
				.b2(W2G028),
				.b3(W2G108),
				.b4(W2G118),
				.b5(W2G128),
				.b6(W2G208),
				.b7(W2G218),
				.b8(W2G228),
				.c(c2812G)
);

ninexnine_unit ninexnine_unit_5357(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2G009),
				.b1(W2G019),
				.b2(W2G029),
				.b3(W2G109),
				.b4(W2G119),
				.b5(W2G129),
				.b6(W2G209),
				.b7(W2G219),
				.b8(W2G229),
				.c(c2912G)
);

ninexnine_unit ninexnine_unit_5358(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2G00A),
				.b1(W2G01A),
				.b2(W2G02A),
				.b3(W2G10A),
				.b4(W2G11A),
				.b5(W2G12A),
				.b6(W2G20A),
				.b7(W2G21A),
				.b8(W2G22A),
				.c(c2A12G)
);

ninexnine_unit ninexnine_unit_5359(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2G00B),
				.b1(W2G01B),
				.b2(W2G02B),
				.b3(W2G10B),
				.b4(W2G11B),
				.b5(W2G12B),
				.b6(W2G20B),
				.b7(W2G21B),
				.b8(W2G22B),
				.c(c2B12G)
);

ninexnine_unit ninexnine_unit_5360(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2G00C),
				.b1(W2G01C),
				.b2(W2G02C),
				.b3(W2G10C),
				.b4(W2G11C),
				.b5(W2G12C),
				.b6(W2G20C),
				.b7(W2G21C),
				.b8(W2G22C),
				.c(c2C12G)
);

ninexnine_unit ninexnine_unit_5361(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2G00D),
				.b1(W2G01D),
				.b2(W2G02D),
				.b3(W2G10D),
				.b4(W2G11D),
				.b5(W2G12D),
				.b6(W2G20D),
				.b7(W2G21D),
				.b8(W2G22D),
				.c(c2D12G)
);

ninexnine_unit ninexnine_unit_5362(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2G00E),
				.b1(W2G01E),
				.b2(W2G02E),
				.b3(W2G10E),
				.b4(W2G11E),
				.b5(W2G12E),
				.b6(W2G20E),
				.b7(W2G21E),
				.b8(W2G22E),
				.c(c2E12G)
);

ninexnine_unit ninexnine_unit_5363(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2G00F),
				.b1(W2G01F),
				.b2(W2G02F),
				.b3(W2G10F),
				.b4(W2G11F),
				.b5(W2G12F),
				.b6(W2G20F),
				.b7(W2G21F),
				.b8(W2G22F),
				.c(c2F12G)
);

assign C212G=c2012G+c2112G+c2212G+c2312G+c2412G+c2512G+c2612G+c2712G+c2812G+c2912G+c2A12G+c2B12G+c2C12G+c2D12G+c2E12G+c2F12G;
assign A212G=(C212G>=0)?1:0;

assign P312G=A212G;

ninexnine_unit ninexnine_unit_5364(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2G000),
				.b1(W2G010),
				.b2(W2G020),
				.b3(W2G100),
				.b4(W2G110),
				.b5(W2G120),
				.b6(W2G200),
				.b7(W2G210),
				.b8(W2G220),
				.c(c2020G)
);

ninexnine_unit ninexnine_unit_5365(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2G001),
				.b1(W2G011),
				.b2(W2G021),
				.b3(W2G101),
				.b4(W2G111),
				.b5(W2G121),
				.b6(W2G201),
				.b7(W2G211),
				.b8(W2G221),
				.c(c2120G)
);

ninexnine_unit ninexnine_unit_5366(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2G002),
				.b1(W2G012),
				.b2(W2G022),
				.b3(W2G102),
				.b4(W2G112),
				.b5(W2G122),
				.b6(W2G202),
				.b7(W2G212),
				.b8(W2G222),
				.c(c2220G)
);

ninexnine_unit ninexnine_unit_5367(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2G003),
				.b1(W2G013),
				.b2(W2G023),
				.b3(W2G103),
				.b4(W2G113),
				.b5(W2G123),
				.b6(W2G203),
				.b7(W2G213),
				.b8(W2G223),
				.c(c2320G)
);

ninexnine_unit ninexnine_unit_5368(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2G004),
				.b1(W2G014),
				.b2(W2G024),
				.b3(W2G104),
				.b4(W2G114),
				.b5(W2G124),
				.b6(W2G204),
				.b7(W2G214),
				.b8(W2G224),
				.c(c2420G)
);

ninexnine_unit ninexnine_unit_5369(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2G005),
				.b1(W2G015),
				.b2(W2G025),
				.b3(W2G105),
				.b4(W2G115),
				.b5(W2G125),
				.b6(W2G205),
				.b7(W2G215),
				.b8(W2G225),
				.c(c2520G)
);

ninexnine_unit ninexnine_unit_5370(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2G006),
				.b1(W2G016),
				.b2(W2G026),
				.b3(W2G106),
				.b4(W2G116),
				.b5(W2G126),
				.b6(W2G206),
				.b7(W2G216),
				.b8(W2G226),
				.c(c2620G)
);

ninexnine_unit ninexnine_unit_5371(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2G007),
				.b1(W2G017),
				.b2(W2G027),
				.b3(W2G107),
				.b4(W2G117),
				.b5(W2G127),
				.b6(W2G207),
				.b7(W2G217),
				.b8(W2G227),
				.c(c2720G)
);

ninexnine_unit ninexnine_unit_5372(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2G008),
				.b1(W2G018),
				.b2(W2G028),
				.b3(W2G108),
				.b4(W2G118),
				.b5(W2G128),
				.b6(W2G208),
				.b7(W2G218),
				.b8(W2G228),
				.c(c2820G)
);

ninexnine_unit ninexnine_unit_5373(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2G009),
				.b1(W2G019),
				.b2(W2G029),
				.b3(W2G109),
				.b4(W2G119),
				.b5(W2G129),
				.b6(W2G209),
				.b7(W2G219),
				.b8(W2G229),
				.c(c2920G)
);

ninexnine_unit ninexnine_unit_5374(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2G00A),
				.b1(W2G01A),
				.b2(W2G02A),
				.b3(W2G10A),
				.b4(W2G11A),
				.b5(W2G12A),
				.b6(W2G20A),
				.b7(W2G21A),
				.b8(W2G22A),
				.c(c2A20G)
);

ninexnine_unit ninexnine_unit_5375(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2G00B),
				.b1(W2G01B),
				.b2(W2G02B),
				.b3(W2G10B),
				.b4(W2G11B),
				.b5(W2G12B),
				.b6(W2G20B),
				.b7(W2G21B),
				.b8(W2G22B),
				.c(c2B20G)
);

ninexnine_unit ninexnine_unit_5376(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2G00C),
				.b1(W2G01C),
				.b2(W2G02C),
				.b3(W2G10C),
				.b4(W2G11C),
				.b5(W2G12C),
				.b6(W2G20C),
				.b7(W2G21C),
				.b8(W2G22C),
				.c(c2C20G)
);

ninexnine_unit ninexnine_unit_5377(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2G00D),
				.b1(W2G01D),
				.b2(W2G02D),
				.b3(W2G10D),
				.b4(W2G11D),
				.b5(W2G12D),
				.b6(W2G20D),
				.b7(W2G21D),
				.b8(W2G22D),
				.c(c2D20G)
);

ninexnine_unit ninexnine_unit_5378(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2G00E),
				.b1(W2G01E),
				.b2(W2G02E),
				.b3(W2G10E),
				.b4(W2G11E),
				.b5(W2G12E),
				.b6(W2G20E),
				.b7(W2G21E),
				.b8(W2G22E),
				.c(c2E20G)
);

ninexnine_unit ninexnine_unit_5379(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2G00F),
				.b1(W2G01F),
				.b2(W2G02F),
				.b3(W2G10F),
				.b4(W2G11F),
				.b5(W2G12F),
				.b6(W2G20F),
				.b7(W2G21F),
				.b8(W2G22F),
				.c(c2F20G)
);

assign C220G=c2020G+c2120G+c2220G+c2320G+c2420G+c2520G+c2620G+c2720G+c2820G+c2920G+c2A20G+c2B20G+c2C20G+c2D20G+c2E20G+c2F20G;
assign A220G=(C220G>=0)?1:0;

assign P320G=A220G;

ninexnine_unit ninexnine_unit_5380(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2G000),
				.b1(W2G010),
				.b2(W2G020),
				.b3(W2G100),
				.b4(W2G110),
				.b5(W2G120),
				.b6(W2G200),
				.b7(W2G210),
				.b8(W2G220),
				.c(c2021G)
);

ninexnine_unit ninexnine_unit_5381(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2G001),
				.b1(W2G011),
				.b2(W2G021),
				.b3(W2G101),
				.b4(W2G111),
				.b5(W2G121),
				.b6(W2G201),
				.b7(W2G211),
				.b8(W2G221),
				.c(c2121G)
);

ninexnine_unit ninexnine_unit_5382(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2G002),
				.b1(W2G012),
				.b2(W2G022),
				.b3(W2G102),
				.b4(W2G112),
				.b5(W2G122),
				.b6(W2G202),
				.b7(W2G212),
				.b8(W2G222),
				.c(c2221G)
);

ninexnine_unit ninexnine_unit_5383(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2G003),
				.b1(W2G013),
				.b2(W2G023),
				.b3(W2G103),
				.b4(W2G113),
				.b5(W2G123),
				.b6(W2G203),
				.b7(W2G213),
				.b8(W2G223),
				.c(c2321G)
);

ninexnine_unit ninexnine_unit_5384(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2G004),
				.b1(W2G014),
				.b2(W2G024),
				.b3(W2G104),
				.b4(W2G114),
				.b5(W2G124),
				.b6(W2G204),
				.b7(W2G214),
				.b8(W2G224),
				.c(c2421G)
);

ninexnine_unit ninexnine_unit_5385(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2G005),
				.b1(W2G015),
				.b2(W2G025),
				.b3(W2G105),
				.b4(W2G115),
				.b5(W2G125),
				.b6(W2G205),
				.b7(W2G215),
				.b8(W2G225),
				.c(c2521G)
);

ninexnine_unit ninexnine_unit_5386(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2G006),
				.b1(W2G016),
				.b2(W2G026),
				.b3(W2G106),
				.b4(W2G116),
				.b5(W2G126),
				.b6(W2G206),
				.b7(W2G216),
				.b8(W2G226),
				.c(c2621G)
);

ninexnine_unit ninexnine_unit_5387(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2G007),
				.b1(W2G017),
				.b2(W2G027),
				.b3(W2G107),
				.b4(W2G117),
				.b5(W2G127),
				.b6(W2G207),
				.b7(W2G217),
				.b8(W2G227),
				.c(c2721G)
);

ninexnine_unit ninexnine_unit_5388(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2G008),
				.b1(W2G018),
				.b2(W2G028),
				.b3(W2G108),
				.b4(W2G118),
				.b5(W2G128),
				.b6(W2G208),
				.b7(W2G218),
				.b8(W2G228),
				.c(c2821G)
);

ninexnine_unit ninexnine_unit_5389(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2G009),
				.b1(W2G019),
				.b2(W2G029),
				.b3(W2G109),
				.b4(W2G119),
				.b5(W2G129),
				.b6(W2G209),
				.b7(W2G219),
				.b8(W2G229),
				.c(c2921G)
);

ninexnine_unit ninexnine_unit_5390(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2G00A),
				.b1(W2G01A),
				.b2(W2G02A),
				.b3(W2G10A),
				.b4(W2G11A),
				.b5(W2G12A),
				.b6(W2G20A),
				.b7(W2G21A),
				.b8(W2G22A),
				.c(c2A21G)
);

ninexnine_unit ninexnine_unit_5391(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2G00B),
				.b1(W2G01B),
				.b2(W2G02B),
				.b3(W2G10B),
				.b4(W2G11B),
				.b5(W2G12B),
				.b6(W2G20B),
				.b7(W2G21B),
				.b8(W2G22B),
				.c(c2B21G)
);

ninexnine_unit ninexnine_unit_5392(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2G00C),
				.b1(W2G01C),
				.b2(W2G02C),
				.b3(W2G10C),
				.b4(W2G11C),
				.b5(W2G12C),
				.b6(W2G20C),
				.b7(W2G21C),
				.b8(W2G22C),
				.c(c2C21G)
);

ninexnine_unit ninexnine_unit_5393(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2G00D),
				.b1(W2G01D),
				.b2(W2G02D),
				.b3(W2G10D),
				.b4(W2G11D),
				.b5(W2G12D),
				.b6(W2G20D),
				.b7(W2G21D),
				.b8(W2G22D),
				.c(c2D21G)
);

ninexnine_unit ninexnine_unit_5394(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2G00E),
				.b1(W2G01E),
				.b2(W2G02E),
				.b3(W2G10E),
				.b4(W2G11E),
				.b5(W2G12E),
				.b6(W2G20E),
				.b7(W2G21E),
				.b8(W2G22E),
				.c(c2E21G)
);

ninexnine_unit ninexnine_unit_5395(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2G00F),
				.b1(W2G01F),
				.b2(W2G02F),
				.b3(W2G10F),
				.b4(W2G11F),
				.b5(W2G12F),
				.b6(W2G20F),
				.b7(W2G21F),
				.b8(W2G22F),
				.c(c2F21G)
);

assign C221G=c2021G+c2121G+c2221G+c2321G+c2421G+c2521G+c2621G+c2721G+c2821G+c2921G+c2A21G+c2B21G+c2C21G+c2D21G+c2E21G+c2F21G;
assign A221G=(C221G>=0)?1:0;

assign P321G=A221G;

ninexnine_unit ninexnine_unit_5396(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2G000),
				.b1(W2G010),
				.b2(W2G020),
				.b3(W2G100),
				.b4(W2G110),
				.b5(W2G120),
				.b6(W2G200),
				.b7(W2G210),
				.b8(W2G220),
				.c(c2022G)
);

ninexnine_unit ninexnine_unit_5397(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2G001),
				.b1(W2G011),
				.b2(W2G021),
				.b3(W2G101),
				.b4(W2G111),
				.b5(W2G121),
				.b6(W2G201),
				.b7(W2G211),
				.b8(W2G221),
				.c(c2122G)
);

ninexnine_unit ninexnine_unit_5398(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2G002),
				.b1(W2G012),
				.b2(W2G022),
				.b3(W2G102),
				.b4(W2G112),
				.b5(W2G122),
				.b6(W2G202),
				.b7(W2G212),
				.b8(W2G222),
				.c(c2222G)
);

ninexnine_unit ninexnine_unit_5399(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2G003),
				.b1(W2G013),
				.b2(W2G023),
				.b3(W2G103),
				.b4(W2G113),
				.b5(W2G123),
				.b6(W2G203),
				.b7(W2G213),
				.b8(W2G223),
				.c(c2322G)
);

ninexnine_unit ninexnine_unit_5400(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2G004),
				.b1(W2G014),
				.b2(W2G024),
				.b3(W2G104),
				.b4(W2G114),
				.b5(W2G124),
				.b6(W2G204),
				.b7(W2G214),
				.b8(W2G224),
				.c(c2422G)
);

ninexnine_unit ninexnine_unit_5401(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2G005),
				.b1(W2G015),
				.b2(W2G025),
				.b3(W2G105),
				.b4(W2G115),
				.b5(W2G125),
				.b6(W2G205),
				.b7(W2G215),
				.b8(W2G225),
				.c(c2522G)
);

ninexnine_unit ninexnine_unit_5402(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2G006),
				.b1(W2G016),
				.b2(W2G026),
				.b3(W2G106),
				.b4(W2G116),
				.b5(W2G126),
				.b6(W2G206),
				.b7(W2G216),
				.b8(W2G226),
				.c(c2622G)
);

ninexnine_unit ninexnine_unit_5403(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2G007),
				.b1(W2G017),
				.b2(W2G027),
				.b3(W2G107),
				.b4(W2G117),
				.b5(W2G127),
				.b6(W2G207),
				.b7(W2G217),
				.b8(W2G227),
				.c(c2722G)
);

ninexnine_unit ninexnine_unit_5404(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2G008),
				.b1(W2G018),
				.b2(W2G028),
				.b3(W2G108),
				.b4(W2G118),
				.b5(W2G128),
				.b6(W2G208),
				.b7(W2G218),
				.b8(W2G228),
				.c(c2822G)
);

ninexnine_unit ninexnine_unit_5405(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2G009),
				.b1(W2G019),
				.b2(W2G029),
				.b3(W2G109),
				.b4(W2G119),
				.b5(W2G129),
				.b6(W2G209),
				.b7(W2G219),
				.b8(W2G229),
				.c(c2922G)
);

ninexnine_unit ninexnine_unit_5406(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2G00A),
				.b1(W2G01A),
				.b2(W2G02A),
				.b3(W2G10A),
				.b4(W2G11A),
				.b5(W2G12A),
				.b6(W2G20A),
				.b7(W2G21A),
				.b8(W2G22A),
				.c(c2A22G)
);

ninexnine_unit ninexnine_unit_5407(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2G00B),
				.b1(W2G01B),
				.b2(W2G02B),
				.b3(W2G10B),
				.b4(W2G11B),
				.b5(W2G12B),
				.b6(W2G20B),
				.b7(W2G21B),
				.b8(W2G22B),
				.c(c2B22G)
);

ninexnine_unit ninexnine_unit_5408(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2G00C),
				.b1(W2G01C),
				.b2(W2G02C),
				.b3(W2G10C),
				.b4(W2G11C),
				.b5(W2G12C),
				.b6(W2G20C),
				.b7(W2G21C),
				.b8(W2G22C),
				.c(c2C22G)
);

ninexnine_unit ninexnine_unit_5409(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2G00D),
				.b1(W2G01D),
				.b2(W2G02D),
				.b3(W2G10D),
				.b4(W2G11D),
				.b5(W2G12D),
				.b6(W2G20D),
				.b7(W2G21D),
				.b8(W2G22D),
				.c(c2D22G)
);

ninexnine_unit ninexnine_unit_5410(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2G00E),
				.b1(W2G01E),
				.b2(W2G02E),
				.b3(W2G10E),
				.b4(W2G11E),
				.b5(W2G12E),
				.b6(W2G20E),
				.b7(W2G21E),
				.b8(W2G22E),
				.c(c2E22G)
);

ninexnine_unit ninexnine_unit_5411(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2G00F),
				.b1(W2G01F),
				.b2(W2G02F),
				.b3(W2G10F),
				.b4(W2G11F),
				.b5(W2G12F),
				.b6(W2G20F),
				.b7(W2G21F),
				.b8(W2G22F),
				.c(c2F22G)
);

assign C222G=c2022G+c2122G+c2222G+c2322G+c2422G+c2522G+c2622G+c2722G+c2822G+c2922G+c2A22G+c2B22G+c2C22G+c2D22G+c2E22G+c2F22G;
assign A222G=(C222G>=0)?1:0;

assign P322G=A222G;

ninexnine_unit ninexnine_unit_5412(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2H000),
				.b1(W2H010),
				.b2(W2H020),
				.b3(W2H100),
				.b4(W2H110),
				.b5(W2H120),
				.b6(W2H200),
				.b7(W2H210),
				.b8(W2H220),
				.c(c2000H)
);

ninexnine_unit ninexnine_unit_5413(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2H001),
				.b1(W2H011),
				.b2(W2H021),
				.b3(W2H101),
				.b4(W2H111),
				.b5(W2H121),
				.b6(W2H201),
				.b7(W2H211),
				.b8(W2H221),
				.c(c2100H)
);

ninexnine_unit ninexnine_unit_5414(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2H002),
				.b1(W2H012),
				.b2(W2H022),
				.b3(W2H102),
				.b4(W2H112),
				.b5(W2H122),
				.b6(W2H202),
				.b7(W2H212),
				.b8(W2H222),
				.c(c2200H)
);

ninexnine_unit ninexnine_unit_5415(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2H003),
				.b1(W2H013),
				.b2(W2H023),
				.b3(W2H103),
				.b4(W2H113),
				.b5(W2H123),
				.b6(W2H203),
				.b7(W2H213),
				.b8(W2H223),
				.c(c2300H)
);

ninexnine_unit ninexnine_unit_5416(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2H004),
				.b1(W2H014),
				.b2(W2H024),
				.b3(W2H104),
				.b4(W2H114),
				.b5(W2H124),
				.b6(W2H204),
				.b7(W2H214),
				.b8(W2H224),
				.c(c2400H)
);

ninexnine_unit ninexnine_unit_5417(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2H005),
				.b1(W2H015),
				.b2(W2H025),
				.b3(W2H105),
				.b4(W2H115),
				.b5(W2H125),
				.b6(W2H205),
				.b7(W2H215),
				.b8(W2H225),
				.c(c2500H)
);

ninexnine_unit ninexnine_unit_5418(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2H006),
				.b1(W2H016),
				.b2(W2H026),
				.b3(W2H106),
				.b4(W2H116),
				.b5(W2H126),
				.b6(W2H206),
				.b7(W2H216),
				.b8(W2H226),
				.c(c2600H)
);

ninexnine_unit ninexnine_unit_5419(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2H007),
				.b1(W2H017),
				.b2(W2H027),
				.b3(W2H107),
				.b4(W2H117),
				.b5(W2H127),
				.b6(W2H207),
				.b7(W2H217),
				.b8(W2H227),
				.c(c2700H)
);

ninexnine_unit ninexnine_unit_5420(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2H008),
				.b1(W2H018),
				.b2(W2H028),
				.b3(W2H108),
				.b4(W2H118),
				.b5(W2H128),
				.b6(W2H208),
				.b7(W2H218),
				.b8(W2H228),
				.c(c2800H)
);

ninexnine_unit ninexnine_unit_5421(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2H009),
				.b1(W2H019),
				.b2(W2H029),
				.b3(W2H109),
				.b4(W2H119),
				.b5(W2H129),
				.b6(W2H209),
				.b7(W2H219),
				.b8(W2H229),
				.c(c2900H)
);

ninexnine_unit ninexnine_unit_5422(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2H00A),
				.b1(W2H01A),
				.b2(W2H02A),
				.b3(W2H10A),
				.b4(W2H11A),
				.b5(W2H12A),
				.b6(W2H20A),
				.b7(W2H21A),
				.b8(W2H22A),
				.c(c2A00H)
);

ninexnine_unit ninexnine_unit_5423(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2H00B),
				.b1(W2H01B),
				.b2(W2H02B),
				.b3(W2H10B),
				.b4(W2H11B),
				.b5(W2H12B),
				.b6(W2H20B),
				.b7(W2H21B),
				.b8(W2H22B),
				.c(c2B00H)
);

ninexnine_unit ninexnine_unit_5424(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2H00C),
				.b1(W2H01C),
				.b2(W2H02C),
				.b3(W2H10C),
				.b4(W2H11C),
				.b5(W2H12C),
				.b6(W2H20C),
				.b7(W2H21C),
				.b8(W2H22C),
				.c(c2C00H)
);

ninexnine_unit ninexnine_unit_5425(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2H00D),
				.b1(W2H01D),
				.b2(W2H02D),
				.b3(W2H10D),
				.b4(W2H11D),
				.b5(W2H12D),
				.b6(W2H20D),
				.b7(W2H21D),
				.b8(W2H22D),
				.c(c2D00H)
);

ninexnine_unit ninexnine_unit_5426(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2H00E),
				.b1(W2H01E),
				.b2(W2H02E),
				.b3(W2H10E),
				.b4(W2H11E),
				.b5(W2H12E),
				.b6(W2H20E),
				.b7(W2H21E),
				.b8(W2H22E),
				.c(c2E00H)
);

ninexnine_unit ninexnine_unit_5427(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2H00F),
				.b1(W2H01F),
				.b2(W2H02F),
				.b3(W2H10F),
				.b4(W2H11F),
				.b5(W2H12F),
				.b6(W2H20F),
				.b7(W2H21F),
				.b8(W2H22F),
				.c(c2F00H)
);

assign C200H=c2000H+c2100H+c2200H+c2300H+c2400H+c2500H+c2600H+c2700H+c2800H+c2900H+c2A00H+c2B00H+c2C00H+c2D00H+c2E00H+c2F00H;
assign A200H=(C200H>=0)?1:0;

assign P300H=A200H;

ninexnine_unit ninexnine_unit_5428(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2H000),
				.b1(W2H010),
				.b2(W2H020),
				.b3(W2H100),
				.b4(W2H110),
				.b5(W2H120),
				.b6(W2H200),
				.b7(W2H210),
				.b8(W2H220),
				.c(c2001H)
);

ninexnine_unit ninexnine_unit_5429(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2H001),
				.b1(W2H011),
				.b2(W2H021),
				.b3(W2H101),
				.b4(W2H111),
				.b5(W2H121),
				.b6(W2H201),
				.b7(W2H211),
				.b8(W2H221),
				.c(c2101H)
);

ninexnine_unit ninexnine_unit_5430(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2H002),
				.b1(W2H012),
				.b2(W2H022),
				.b3(W2H102),
				.b4(W2H112),
				.b5(W2H122),
				.b6(W2H202),
				.b7(W2H212),
				.b8(W2H222),
				.c(c2201H)
);

ninexnine_unit ninexnine_unit_5431(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2H003),
				.b1(W2H013),
				.b2(W2H023),
				.b3(W2H103),
				.b4(W2H113),
				.b5(W2H123),
				.b6(W2H203),
				.b7(W2H213),
				.b8(W2H223),
				.c(c2301H)
);

ninexnine_unit ninexnine_unit_5432(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2H004),
				.b1(W2H014),
				.b2(W2H024),
				.b3(W2H104),
				.b4(W2H114),
				.b5(W2H124),
				.b6(W2H204),
				.b7(W2H214),
				.b8(W2H224),
				.c(c2401H)
);

ninexnine_unit ninexnine_unit_5433(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2H005),
				.b1(W2H015),
				.b2(W2H025),
				.b3(W2H105),
				.b4(W2H115),
				.b5(W2H125),
				.b6(W2H205),
				.b7(W2H215),
				.b8(W2H225),
				.c(c2501H)
);

ninexnine_unit ninexnine_unit_5434(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2H006),
				.b1(W2H016),
				.b2(W2H026),
				.b3(W2H106),
				.b4(W2H116),
				.b5(W2H126),
				.b6(W2H206),
				.b7(W2H216),
				.b8(W2H226),
				.c(c2601H)
);

ninexnine_unit ninexnine_unit_5435(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2H007),
				.b1(W2H017),
				.b2(W2H027),
				.b3(W2H107),
				.b4(W2H117),
				.b5(W2H127),
				.b6(W2H207),
				.b7(W2H217),
				.b8(W2H227),
				.c(c2701H)
);

ninexnine_unit ninexnine_unit_5436(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2H008),
				.b1(W2H018),
				.b2(W2H028),
				.b3(W2H108),
				.b4(W2H118),
				.b5(W2H128),
				.b6(W2H208),
				.b7(W2H218),
				.b8(W2H228),
				.c(c2801H)
);

ninexnine_unit ninexnine_unit_5437(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2H009),
				.b1(W2H019),
				.b2(W2H029),
				.b3(W2H109),
				.b4(W2H119),
				.b5(W2H129),
				.b6(W2H209),
				.b7(W2H219),
				.b8(W2H229),
				.c(c2901H)
);

ninexnine_unit ninexnine_unit_5438(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2H00A),
				.b1(W2H01A),
				.b2(W2H02A),
				.b3(W2H10A),
				.b4(W2H11A),
				.b5(W2H12A),
				.b6(W2H20A),
				.b7(W2H21A),
				.b8(W2H22A),
				.c(c2A01H)
);

ninexnine_unit ninexnine_unit_5439(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2H00B),
				.b1(W2H01B),
				.b2(W2H02B),
				.b3(W2H10B),
				.b4(W2H11B),
				.b5(W2H12B),
				.b6(W2H20B),
				.b7(W2H21B),
				.b8(W2H22B),
				.c(c2B01H)
);

ninexnine_unit ninexnine_unit_5440(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2H00C),
				.b1(W2H01C),
				.b2(W2H02C),
				.b3(W2H10C),
				.b4(W2H11C),
				.b5(W2H12C),
				.b6(W2H20C),
				.b7(W2H21C),
				.b8(W2H22C),
				.c(c2C01H)
);

ninexnine_unit ninexnine_unit_5441(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2H00D),
				.b1(W2H01D),
				.b2(W2H02D),
				.b3(W2H10D),
				.b4(W2H11D),
				.b5(W2H12D),
				.b6(W2H20D),
				.b7(W2H21D),
				.b8(W2H22D),
				.c(c2D01H)
);

ninexnine_unit ninexnine_unit_5442(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2H00E),
				.b1(W2H01E),
				.b2(W2H02E),
				.b3(W2H10E),
				.b4(W2H11E),
				.b5(W2H12E),
				.b6(W2H20E),
				.b7(W2H21E),
				.b8(W2H22E),
				.c(c2E01H)
);

ninexnine_unit ninexnine_unit_5443(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2H00F),
				.b1(W2H01F),
				.b2(W2H02F),
				.b3(W2H10F),
				.b4(W2H11F),
				.b5(W2H12F),
				.b6(W2H20F),
				.b7(W2H21F),
				.b8(W2H22F),
				.c(c2F01H)
);

assign C201H=c2001H+c2101H+c2201H+c2301H+c2401H+c2501H+c2601H+c2701H+c2801H+c2901H+c2A01H+c2B01H+c2C01H+c2D01H+c2E01H+c2F01H;
assign A201H=(C201H>=0)?1:0;

assign P301H=A201H;

ninexnine_unit ninexnine_unit_5444(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2H000),
				.b1(W2H010),
				.b2(W2H020),
				.b3(W2H100),
				.b4(W2H110),
				.b5(W2H120),
				.b6(W2H200),
				.b7(W2H210),
				.b8(W2H220),
				.c(c2002H)
);

ninexnine_unit ninexnine_unit_5445(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2H001),
				.b1(W2H011),
				.b2(W2H021),
				.b3(W2H101),
				.b4(W2H111),
				.b5(W2H121),
				.b6(W2H201),
				.b7(W2H211),
				.b8(W2H221),
				.c(c2102H)
);

ninexnine_unit ninexnine_unit_5446(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2H002),
				.b1(W2H012),
				.b2(W2H022),
				.b3(W2H102),
				.b4(W2H112),
				.b5(W2H122),
				.b6(W2H202),
				.b7(W2H212),
				.b8(W2H222),
				.c(c2202H)
);

ninexnine_unit ninexnine_unit_5447(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2H003),
				.b1(W2H013),
				.b2(W2H023),
				.b3(W2H103),
				.b4(W2H113),
				.b5(W2H123),
				.b6(W2H203),
				.b7(W2H213),
				.b8(W2H223),
				.c(c2302H)
);

ninexnine_unit ninexnine_unit_5448(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2H004),
				.b1(W2H014),
				.b2(W2H024),
				.b3(W2H104),
				.b4(W2H114),
				.b5(W2H124),
				.b6(W2H204),
				.b7(W2H214),
				.b8(W2H224),
				.c(c2402H)
);

ninexnine_unit ninexnine_unit_5449(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2H005),
				.b1(W2H015),
				.b2(W2H025),
				.b3(W2H105),
				.b4(W2H115),
				.b5(W2H125),
				.b6(W2H205),
				.b7(W2H215),
				.b8(W2H225),
				.c(c2502H)
);

ninexnine_unit ninexnine_unit_5450(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2H006),
				.b1(W2H016),
				.b2(W2H026),
				.b3(W2H106),
				.b4(W2H116),
				.b5(W2H126),
				.b6(W2H206),
				.b7(W2H216),
				.b8(W2H226),
				.c(c2602H)
);

ninexnine_unit ninexnine_unit_5451(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2H007),
				.b1(W2H017),
				.b2(W2H027),
				.b3(W2H107),
				.b4(W2H117),
				.b5(W2H127),
				.b6(W2H207),
				.b7(W2H217),
				.b8(W2H227),
				.c(c2702H)
);

ninexnine_unit ninexnine_unit_5452(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2H008),
				.b1(W2H018),
				.b2(W2H028),
				.b3(W2H108),
				.b4(W2H118),
				.b5(W2H128),
				.b6(W2H208),
				.b7(W2H218),
				.b8(W2H228),
				.c(c2802H)
);

ninexnine_unit ninexnine_unit_5453(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2H009),
				.b1(W2H019),
				.b2(W2H029),
				.b3(W2H109),
				.b4(W2H119),
				.b5(W2H129),
				.b6(W2H209),
				.b7(W2H219),
				.b8(W2H229),
				.c(c2902H)
);

ninexnine_unit ninexnine_unit_5454(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2H00A),
				.b1(W2H01A),
				.b2(W2H02A),
				.b3(W2H10A),
				.b4(W2H11A),
				.b5(W2H12A),
				.b6(W2H20A),
				.b7(W2H21A),
				.b8(W2H22A),
				.c(c2A02H)
);

ninexnine_unit ninexnine_unit_5455(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2H00B),
				.b1(W2H01B),
				.b2(W2H02B),
				.b3(W2H10B),
				.b4(W2H11B),
				.b5(W2H12B),
				.b6(W2H20B),
				.b7(W2H21B),
				.b8(W2H22B),
				.c(c2B02H)
);

ninexnine_unit ninexnine_unit_5456(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2H00C),
				.b1(W2H01C),
				.b2(W2H02C),
				.b3(W2H10C),
				.b4(W2H11C),
				.b5(W2H12C),
				.b6(W2H20C),
				.b7(W2H21C),
				.b8(W2H22C),
				.c(c2C02H)
);

ninexnine_unit ninexnine_unit_5457(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2H00D),
				.b1(W2H01D),
				.b2(W2H02D),
				.b3(W2H10D),
				.b4(W2H11D),
				.b5(W2H12D),
				.b6(W2H20D),
				.b7(W2H21D),
				.b8(W2H22D),
				.c(c2D02H)
);

ninexnine_unit ninexnine_unit_5458(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2H00E),
				.b1(W2H01E),
				.b2(W2H02E),
				.b3(W2H10E),
				.b4(W2H11E),
				.b5(W2H12E),
				.b6(W2H20E),
				.b7(W2H21E),
				.b8(W2H22E),
				.c(c2E02H)
);

ninexnine_unit ninexnine_unit_5459(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2H00F),
				.b1(W2H01F),
				.b2(W2H02F),
				.b3(W2H10F),
				.b4(W2H11F),
				.b5(W2H12F),
				.b6(W2H20F),
				.b7(W2H21F),
				.b8(W2H22F),
				.c(c2F02H)
);

assign C202H=c2002H+c2102H+c2202H+c2302H+c2402H+c2502H+c2602H+c2702H+c2802H+c2902H+c2A02H+c2B02H+c2C02H+c2D02H+c2E02H+c2F02H;
assign A202H=(C202H>=0)?1:0;

assign P302H=A202H;

ninexnine_unit ninexnine_unit_5460(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2H000),
				.b1(W2H010),
				.b2(W2H020),
				.b3(W2H100),
				.b4(W2H110),
				.b5(W2H120),
				.b6(W2H200),
				.b7(W2H210),
				.b8(W2H220),
				.c(c2010H)
);

ninexnine_unit ninexnine_unit_5461(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2H001),
				.b1(W2H011),
				.b2(W2H021),
				.b3(W2H101),
				.b4(W2H111),
				.b5(W2H121),
				.b6(W2H201),
				.b7(W2H211),
				.b8(W2H221),
				.c(c2110H)
);

ninexnine_unit ninexnine_unit_5462(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2H002),
				.b1(W2H012),
				.b2(W2H022),
				.b3(W2H102),
				.b4(W2H112),
				.b5(W2H122),
				.b6(W2H202),
				.b7(W2H212),
				.b8(W2H222),
				.c(c2210H)
);

ninexnine_unit ninexnine_unit_5463(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2H003),
				.b1(W2H013),
				.b2(W2H023),
				.b3(W2H103),
				.b4(W2H113),
				.b5(W2H123),
				.b6(W2H203),
				.b7(W2H213),
				.b8(W2H223),
				.c(c2310H)
);

ninexnine_unit ninexnine_unit_5464(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2H004),
				.b1(W2H014),
				.b2(W2H024),
				.b3(W2H104),
				.b4(W2H114),
				.b5(W2H124),
				.b6(W2H204),
				.b7(W2H214),
				.b8(W2H224),
				.c(c2410H)
);

ninexnine_unit ninexnine_unit_5465(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2H005),
				.b1(W2H015),
				.b2(W2H025),
				.b3(W2H105),
				.b4(W2H115),
				.b5(W2H125),
				.b6(W2H205),
				.b7(W2H215),
				.b8(W2H225),
				.c(c2510H)
);

ninexnine_unit ninexnine_unit_5466(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2H006),
				.b1(W2H016),
				.b2(W2H026),
				.b3(W2H106),
				.b4(W2H116),
				.b5(W2H126),
				.b6(W2H206),
				.b7(W2H216),
				.b8(W2H226),
				.c(c2610H)
);

ninexnine_unit ninexnine_unit_5467(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2H007),
				.b1(W2H017),
				.b2(W2H027),
				.b3(W2H107),
				.b4(W2H117),
				.b5(W2H127),
				.b6(W2H207),
				.b7(W2H217),
				.b8(W2H227),
				.c(c2710H)
);

ninexnine_unit ninexnine_unit_5468(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2H008),
				.b1(W2H018),
				.b2(W2H028),
				.b3(W2H108),
				.b4(W2H118),
				.b5(W2H128),
				.b6(W2H208),
				.b7(W2H218),
				.b8(W2H228),
				.c(c2810H)
);

ninexnine_unit ninexnine_unit_5469(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2H009),
				.b1(W2H019),
				.b2(W2H029),
				.b3(W2H109),
				.b4(W2H119),
				.b5(W2H129),
				.b6(W2H209),
				.b7(W2H219),
				.b8(W2H229),
				.c(c2910H)
);

ninexnine_unit ninexnine_unit_5470(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2H00A),
				.b1(W2H01A),
				.b2(W2H02A),
				.b3(W2H10A),
				.b4(W2H11A),
				.b5(W2H12A),
				.b6(W2H20A),
				.b7(W2H21A),
				.b8(W2H22A),
				.c(c2A10H)
);

ninexnine_unit ninexnine_unit_5471(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2H00B),
				.b1(W2H01B),
				.b2(W2H02B),
				.b3(W2H10B),
				.b4(W2H11B),
				.b5(W2H12B),
				.b6(W2H20B),
				.b7(W2H21B),
				.b8(W2H22B),
				.c(c2B10H)
);

ninexnine_unit ninexnine_unit_5472(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2H00C),
				.b1(W2H01C),
				.b2(W2H02C),
				.b3(W2H10C),
				.b4(W2H11C),
				.b5(W2H12C),
				.b6(W2H20C),
				.b7(W2H21C),
				.b8(W2H22C),
				.c(c2C10H)
);

ninexnine_unit ninexnine_unit_5473(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2H00D),
				.b1(W2H01D),
				.b2(W2H02D),
				.b3(W2H10D),
				.b4(W2H11D),
				.b5(W2H12D),
				.b6(W2H20D),
				.b7(W2H21D),
				.b8(W2H22D),
				.c(c2D10H)
);

ninexnine_unit ninexnine_unit_5474(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2H00E),
				.b1(W2H01E),
				.b2(W2H02E),
				.b3(W2H10E),
				.b4(W2H11E),
				.b5(W2H12E),
				.b6(W2H20E),
				.b7(W2H21E),
				.b8(W2H22E),
				.c(c2E10H)
);

ninexnine_unit ninexnine_unit_5475(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2H00F),
				.b1(W2H01F),
				.b2(W2H02F),
				.b3(W2H10F),
				.b4(W2H11F),
				.b5(W2H12F),
				.b6(W2H20F),
				.b7(W2H21F),
				.b8(W2H22F),
				.c(c2F10H)
);

assign C210H=c2010H+c2110H+c2210H+c2310H+c2410H+c2510H+c2610H+c2710H+c2810H+c2910H+c2A10H+c2B10H+c2C10H+c2D10H+c2E10H+c2F10H;
assign A210H=(C210H>=0)?1:0;

assign P310H=A210H;

ninexnine_unit ninexnine_unit_5476(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2H000),
				.b1(W2H010),
				.b2(W2H020),
				.b3(W2H100),
				.b4(W2H110),
				.b5(W2H120),
				.b6(W2H200),
				.b7(W2H210),
				.b8(W2H220),
				.c(c2011H)
);

ninexnine_unit ninexnine_unit_5477(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2H001),
				.b1(W2H011),
				.b2(W2H021),
				.b3(W2H101),
				.b4(W2H111),
				.b5(W2H121),
				.b6(W2H201),
				.b7(W2H211),
				.b8(W2H221),
				.c(c2111H)
);

ninexnine_unit ninexnine_unit_5478(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2H002),
				.b1(W2H012),
				.b2(W2H022),
				.b3(W2H102),
				.b4(W2H112),
				.b5(W2H122),
				.b6(W2H202),
				.b7(W2H212),
				.b8(W2H222),
				.c(c2211H)
);

ninexnine_unit ninexnine_unit_5479(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2H003),
				.b1(W2H013),
				.b2(W2H023),
				.b3(W2H103),
				.b4(W2H113),
				.b5(W2H123),
				.b6(W2H203),
				.b7(W2H213),
				.b8(W2H223),
				.c(c2311H)
);

ninexnine_unit ninexnine_unit_5480(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2H004),
				.b1(W2H014),
				.b2(W2H024),
				.b3(W2H104),
				.b4(W2H114),
				.b5(W2H124),
				.b6(W2H204),
				.b7(W2H214),
				.b8(W2H224),
				.c(c2411H)
);

ninexnine_unit ninexnine_unit_5481(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2H005),
				.b1(W2H015),
				.b2(W2H025),
				.b3(W2H105),
				.b4(W2H115),
				.b5(W2H125),
				.b6(W2H205),
				.b7(W2H215),
				.b8(W2H225),
				.c(c2511H)
);

ninexnine_unit ninexnine_unit_5482(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2H006),
				.b1(W2H016),
				.b2(W2H026),
				.b3(W2H106),
				.b4(W2H116),
				.b5(W2H126),
				.b6(W2H206),
				.b7(W2H216),
				.b8(W2H226),
				.c(c2611H)
);

ninexnine_unit ninexnine_unit_5483(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2H007),
				.b1(W2H017),
				.b2(W2H027),
				.b3(W2H107),
				.b4(W2H117),
				.b5(W2H127),
				.b6(W2H207),
				.b7(W2H217),
				.b8(W2H227),
				.c(c2711H)
);

ninexnine_unit ninexnine_unit_5484(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2H008),
				.b1(W2H018),
				.b2(W2H028),
				.b3(W2H108),
				.b4(W2H118),
				.b5(W2H128),
				.b6(W2H208),
				.b7(W2H218),
				.b8(W2H228),
				.c(c2811H)
);

ninexnine_unit ninexnine_unit_5485(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2H009),
				.b1(W2H019),
				.b2(W2H029),
				.b3(W2H109),
				.b4(W2H119),
				.b5(W2H129),
				.b6(W2H209),
				.b7(W2H219),
				.b8(W2H229),
				.c(c2911H)
);

ninexnine_unit ninexnine_unit_5486(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2H00A),
				.b1(W2H01A),
				.b2(W2H02A),
				.b3(W2H10A),
				.b4(W2H11A),
				.b5(W2H12A),
				.b6(W2H20A),
				.b7(W2H21A),
				.b8(W2H22A),
				.c(c2A11H)
);

ninexnine_unit ninexnine_unit_5487(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2H00B),
				.b1(W2H01B),
				.b2(W2H02B),
				.b3(W2H10B),
				.b4(W2H11B),
				.b5(W2H12B),
				.b6(W2H20B),
				.b7(W2H21B),
				.b8(W2H22B),
				.c(c2B11H)
);

ninexnine_unit ninexnine_unit_5488(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2H00C),
				.b1(W2H01C),
				.b2(W2H02C),
				.b3(W2H10C),
				.b4(W2H11C),
				.b5(W2H12C),
				.b6(W2H20C),
				.b7(W2H21C),
				.b8(W2H22C),
				.c(c2C11H)
);

ninexnine_unit ninexnine_unit_5489(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2H00D),
				.b1(W2H01D),
				.b2(W2H02D),
				.b3(W2H10D),
				.b4(W2H11D),
				.b5(W2H12D),
				.b6(W2H20D),
				.b7(W2H21D),
				.b8(W2H22D),
				.c(c2D11H)
);

ninexnine_unit ninexnine_unit_5490(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2H00E),
				.b1(W2H01E),
				.b2(W2H02E),
				.b3(W2H10E),
				.b4(W2H11E),
				.b5(W2H12E),
				.b6(W2H20E),
				.b7(W2H21E),
				.b8(W2H22E),
				.c(c2E11H)
);

ninexnine_unit ninexnine_unit_5491(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2H00F),
				.b1(W2H01F),
				.b2(W2H02F),
				.b3(W2H10F),
				.b4(W2H11F),
				.b5(W2H12F),
				.b6(W2H20F),
				.b7(W2H21F),
				.b8(W2H22F),
				.c(c2F11H)
);

assign C211H=c2011H+c2111H+c2211H+c2311H+c2411H+c2511H+c2611H+c2711H+c2811H+c2911H+c2A11H+c2B11H+c2C11H+c2D11H+c2E11H+c2F11H;
assign A211H=(C211H>=0)?1:0;

assign P311H=A211H;

ninexnine_unit ninexnine_unit_5492(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2H000),
				.b1(W2H010),
				.b2(W2H020),
				.b3(W2H100),
				.b4(W2H110),
				.b5(W2H120),
				.b6(W2H200),
				.b7(W2H210),
				.b8(W2H220),
				.c(c2012H)
);

ninexnine_unit ninexnine_unit_5493(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2H001),
				.b1(W2H011),
				.b2(W2H021),
				.b3(W2H101),
				.b4(W2H111),
				.b5(W2H121),
				.b6(W2H201),
				.b7(W2H211),
				.b8(W2H221),
				.c(c2112H)
);

ninexnine_unit ninexnine_unit_5494(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2H002),
				.b1(W2H012),
				.b2(W2H022),
				.b3(W2H102),
				.b4(W2H112),
				.b5(W2H122),
				.b6(W2H202),
				.b7(W2H212),
				.b8(W2H222),
				.c(c2212H)
);

ninexnine_unit ninexnine_unit_5495(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2H003),
				.b1(W2H013),
				.b2(W2H023),
				.b3(W2H103),
				.b4(W2H113),
				.b5(W2H123),
				.b6(W2H203),
				.b7(W2H213),
				.b8(W2H223),
				.c(c2312H)
);

ninexnine_unit ninexnine_unit_5496(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2H004),
				.b1(W2H014),
				.b2(W2H024),
				.b3(W2H104),
				.b4(W2H114),
				.b5(W2H124),
				.b6(W2H204),
				.b7(W2H214),
				.b8(W2H224),
				.c(c2412H)
);

ninexnine_unit ninexnine_unit_5497(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2H005),
				.b1(W2H015),
				.b2(W2H025),
				.b3(W2H105),
				.b4(W2H115),
				.b5(W2H125),
				.b6(W2H205),
				.b7(W2H215),
				.b8(W2H225),
				.c(c2512H)
);

ninexnine_unit ninexnine_unit_5498(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2H006),
				.b1(W2H016),
				.b2(W2H026),
				.b3(W2H106),
				.b4(W2H116),
				.b5(W2H126),
				.b6(W2H206),
				.b7(W2H216),
				.b8(W2H226),
				.c(c2612H)
);

ninexnine_unit ninexnine_unit_5499(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2H007),
				.b1(W2H017),
				.b2(W2H027),
				.b3(W2H107),
				.b4(W2H117),
				.b5(W2H127),
				.b6(W2H207),
				.b7(W2H217),
				.b8(W2H227),
				.c(c2712H)
);

ninexnine_unit ninexnine_unit_5500(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2H008),
				.b1(W2H018),
				.b2(W2H028),
				.b3(W2H108),
				.b4(W2H118),
				.b5(W2H128),
				.b6(W2H208),
				.b7(W2H218),
				.b8(W2H228),
				.c(c2812H)
);

ninexnine_unit ninexnine_unit_5501(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2H009),
				.b1(W2H019),
				.b2(W2H029),
				.b3(W2H109),
				.b4(W2H119),
				.b5(W2H129),
				.b6(W2H209),
				.b7(W2H219),
				.b8(W2H229),
				.c(c2912H)
);

ninexnine_unit ninexnine_unit_5502(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2H00A),
				.b1(W2H01A),
				.b2(W2H02A),
				.b3(W2H10A),
				.b4(W2H11A),
				.b5(W2H12A),
				.b6(W2H20A),
				.b7(W2H21A),
				.b8(W2H22A),
				.c(c2A12H)
);

ninexnine_unit ninexnine_unit_5503(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2H00B),
				.b1(W2H01B),
				.b2(W2H02B),
				.b3(W2H10B),
				.b4(W2H11B),
				.b5(W2H12B),
				.b6(W2H20B),
				.b7(W2H21B),
				.b8(W2H22B),
				.c(c2B12H)
);

ninexnine_unit ninexnine_unit_5504(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2H00C),
				.b1(W2H01C),
				.b2(W2H02C),
				.b3(W2H10C),
				.b4(W2H11C),
				.b5(W2H12C),
				.b6(W2H20C),
				.b7(W2H21C),
				.b8(W2H22C),
				.c(c2C12H)
);

ninexnine_unit ninexnine_unit_5505(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2H00D),
				.b1(W2H01D),
				.b2(W2H02D),
				.b3(W2H10D),
				.b4(W2H11D),
				.b5(W2H12D),
				.b6(W2H20D),
				.b7(W2H21D),
				.b8(W2H22D),
				.c(c2D12H)
);

ninexnine_unit ninexnine_unit_5506(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2H00E),
				.b1(W2H01E),
				.b2(W2H02E),
				.b3(W2H10E),
				.b4(W2H11E),
				.b5(W2H12E),
				.b6(W2H20E),
				.b7(W2H21E),
				.b8(W2H22E),
				.c(c2E12H)
);

ninexnine_unit ninexnine_unit_5507(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2H00F),
				.b1(W2H01F),
				.b2(W2H02F),
				.b3(W2H10F),
				.b4(W2H11F),
				.b5(W2H12F),
				.b6(W2H20F),
				.b7(W2H21F),
				.b8(W2H22F),
				.c(c2F12H)
);

assign C212H=c2012H+c2112H+c2212H+c2312H+c2412H+c2512H+c2612H+c2712H+c2812H+c2912H+c2A12H+c2B12H+c2C12H+c2D12H+c2E12H+c2F12H;
assign A212H=(C212H>=0)?1:0;

assign P312H=A212H;

ninexnine_unit ninexnine_unit_5508(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2H000),
				.b1(W2H010),
				.b2(W2H020),
				.b3(W2H100),
				.b4(W2H110),
				.b5(W2H120),
				.b6(W2H200),
				.b7(W2H210),
				.b8(W2H220),
				.c(c2020H)
);

ninexnine_unit ninexnine_unit_5509(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2H001),
				.b1(W2H011),
				.b2(W2H021),
				.b3(W2H101),
				.b4(W2H111),
				.b5(W2H121),
				.b6(W2H201),
				.b7(W2H211),
				.b8(W2H221),
				.c(c2120H)
);

ninexnine_unit ninexnine_unit_5510(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2H002),
				.b1(W2H012),
				.b2(W2H022),
				.b3(W2H102),
				.b4(W2H112),
				.b5(W2H122),
				.b6(W2H202),
				.b7(W2H212),
				.b8(W2H222),
				.c(c2220H)
);

ninexnine_unit ninexnine_unit_5511(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2H003),
				.b1(W2H013),
				.b2(W2H023),
				.b3(W2H103),
				.b4(W2H113),
				.b5(W2H123),
				.b6(W2H203),
				.b7(W2H213),
				.b8(W2H223),
				.c(c2320H)
);

ninexnine_unit ninexnine_unit_5512(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2H004),
				.b1(W2H014),
				.b2(W2H024),
				.b3(W2H104),
				.b4(W2H114),
				.b5(W2H124),
				.b6(W2H204),
				.b7(W2H214),
				.b8(W2H224),
				.c(c2420H)
);

ninexnine_unit ninexnine_unit_5513(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2H005),
				.b1(W2H015),
				.b2(W2H025),
				.b3(W2H105),
				.b4(W2H115),
				.b5(W2H125),
				.b6(W2H205),
				.b7(W2H215),
				.b8(W2H225),
				.c(c2520H)
);

ninexnine_unit ninexnine_unit_5514(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2H006),
				.b1(W2H016),
				.b2(W2H026),
				.b3(W2H106),
				.b4(W2H116),
				.b5(W2H126),
				.b6(W2H206),
				.b7(W2H216),
				.b8(W2H226),
				.c(c2620H)
);

ninexnine_unit ninexnine_unit_5515(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2H007),
				.b1(W2H017),
				.b2(W2H027),
				.b3(W2H107),
				.b4(W2H117),
				.b5(W2H127),
				.b6(W2H207),
				.b7(W2H217),
				.b8(W2H227),
				.c(c2720H)
);

ninexnine_unit ninexnine_unit_5516(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2H008),
				.b1(W2H018),
				.b2(W2H028),
				.b3(W2H108),
				.b4(W2H118),
				.b5(W2H128),
				.b6(W2H208),
				.b7(W2H218),
				.b8(W2H228),
				.c(c2820H)
);

ninexnine_unit ninexnine_unit_5517(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2H009),
				.b1(W2H019),
				.b2(W2H029),
				.b3(W2H109),
				.b4(W2H119),
				.b5(W2H129),
				.b6(W2H209),
				.b7(W2H219),
				.b8(W2H229),
				.c(c2920H)
);

ninexnine_unit ninexnine_unit_5518(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2H00A),
				.b1(W2H01A),
				.b2(W2H02A),
				.b3(W2H10A),
				.b4(W2H11A),
				.b5(W2H12A),
				.b6(W2H20A),
				.b7(W2H21A),
				.b8(W2H22A),
				.c(c2A20H)
);

ninexnine_unit ninexnine_unit_5519(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2H00B),
				.b1(W2H01B),
				.b2(W2H02B),
				.b3(W2H10B),
				.b4(W2H11B),
				.b5(W2H12B),
				.b6(W2H20B),
				.b7(W2H21B),
				.b8(W2H22B),
				.c(c2B20H)
);

ninexnine_unit ninexnine_unit_5520(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2H00C),
				.b1(W2H01C),
				.b2(W2H02C),
				.b3(W2H10C),
				.b4(W2H11C),
				.b5(W2H12C),
				.b6(W2H20C),
				.b7(W2H21C),
				.b8(W2H22C),
				.c(c2C20H)
);

ninexnine_unit ninexnine_unit_5521(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2H00D),
				.b1(W2H01D),
				.b2(W2H02D),
				.b3(W2H10D),
				.b4(W2H11D),
				.b5(W2H12D),
				.b6(W2H20D),
				.b7(W2H21D),
				.b8(W2H22D),
				.c(c2D20H)
);

ninexnine_unit ninexnine_unit_5522(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2H00E),
				.b1(W2H01E),
				.b2(W2H02E),
				.b3(W2H10E),
				.b4(W2H11E),
				.b5(W2H12E),
				.b6(W2H20E),
				.b7(W2H21E),
				.b8(W2H22E),
				.c(c2E20H)
);

ninexnine_unit ninexnine_unit_5523(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2H00F),
				.b1(W2H01F),
				.b2(W2H02F),
				.b3(W2H10F),
				.b4(W2H11F),
				.b5(W2H12F),
				.b6(W2H20F),
				.b7(W2H21F),
				.b8(W2H22F),
				.c(c2F20H)
);

assign C220H=c2020H+c2120H+c2220H+c2320H+c2420H+c2520H+c2620H+c2720H+c2820H+c2920H+c2A20H+c2B20H+c2C20H+c2D20H+c2E20H+c2F20H;
assign A220H=(C220H>=0)?1:0;

assign P320H=A220H;

ninexnine_unit ninexnine_unit_5524(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2H000),
				.b1(W2H010),
				.b2(W2H020),
				.b3(W2H100),
				.b4(W2H110),
				.b5(W2H120),
				.b6(W2H200),
				.b7(W2H210),
				.b8(W2H220),
				.c(c2021H)
);

ninexnine_unit ninexnine_unit_5525(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2H001),
				.b1(W2H011),
				.b2(W2H021),
				.b3(W2H101),
				.b4(W2H111),
				.b5(W2H121),
				.b6(W2H201),
				.b7(W2H211),
				.b8(W2H221),
				.c(c2121H)
);

ninexnine_unit ninexnine_unit_5526(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2H002),
				.b1(W2H012),
				.b2(W2H022),
				.b3(W2H102),
				.b4(W2H112),
				.b5(W2H122),
				.b6(W2H202),
				.b7(W2H212),
				.b8(W2H222),
				.c(c2221H)
);

ninexnine_unit ninexnine_unit_5527(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2H003),
				.b1(W2H013),
				.b2(W2H023),
				.b3(W2H103),
				.b4(W2H113),
				.b5(W2H123),
				.b6(W2H203),
				.b7(W2H213),
				.b8(W2H223),
				.c(c2321H)
);

ninexnine_unit ninexnine_unit_5528(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2H004),
				.b1(W2H014),
				.b2(W2H024),
				.b3(W2H104),
				.b4(W2H114),
				.b5(W2H124),
				.b6(W2H204),
				.b7(W2H214),
				.b8(W2H224),
				.c(c2421H)
);

ninexnine_unit ninexnine_unit_5529(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2H005),
				.b1(W2H015),
				.b2(W2H025),
				.b3(W2H105),
				.b4(W2H115),
				.b5(W2H125),
				.b6(W2H205),
				.b7(W2H215),
				.b8(W2H225),
				.c(c2521H)
);

ninexnine_unit ninexnine_unit_5530(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2H006),
				.b1(W2H016),
				.b2(W2H026),
				.b3(W2H106),
				.b4(W2H116),
				.b5(W2H126),
				.b6(W2H206),
				.b7(W2H216),
				.b8(W2H226),
				.c(c2621H)
);

ninexnine_unit ninexnine_unit_5531(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2H007),
				.b1(W2H017),
				.b2(W2H027),
				.b3(W2H107),
				.b4(W2H117),
				.b5(W2H127),
				.b6(W2H207),
				.b7(W2H217),
				.b8(W2H227),
				.c(c2721H)
);

ninexnine_unit ninexnine_unit_5532(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2H008),
				.b1(W2H018),
				.b2(W2H028),
				.b3(W2H108),
				.b4(W2H118),
				.b5(W2H128),
				.b6(W2H208),
				.b7(W2H218),
				.b8(W2H228),
				.c(c2821H)
);

ninexnine_unit ninexnine_unit_5533(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2H009),
				.b1(W2H019),
				.b2(W2H029),
				.b3(W2H109),
				.b4(W2H119),
				.b5(W2H129),
				.b6(W2H209),
				.b7(W2H219),
				.b8(W2H229),
				.c(c2921H)
);

ninexnine_unit ninexnine_unit_5534(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2H00A),
				.b1(W2H01A),
				.b2(W2H02A),
				.b3(W2H10A),
				.b4(W2H11A),
				.b5(W2H12A),
				.b6(W2H20A),
				.b7(W2H21A),
				.b8(W2H22A),
				.c(c2A21H)
);

ninexnine_unit ninexnine_unit_5535(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2H00B),
				.b1(W2H01B),
				.b2(W2H02B),
				.b3(W2H10B),
				.b4(W2H11B),
				.b5(W2H12B),
				.b6(W2H20B),
				.b7(W2H21B),
				.b8(W2H22B),
				.c(c2B21H)
);

ninexnine_unit ninexnine_unit_5536(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2H00C),
				.b1(W2H01C),
				.b2(W2H02C),
				.b3(W2H10C),
				.b4(W2H11C),
				.b5(W2H12C),
				.b6(W2H20C),
				.b7(W2H21C),
				.b8(W2H22C),
				.c(c2C21H)
);

ninexnine_unit ninexnine_unit_5537(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2H00D),
				.b1(W2H01D),
				.b2(W2H02D),
				.b3(W2H10D),
				.b4(W2H11D),
				.b5(W2H12D),
				.b6(W2H20D),
				.b7(W2H21D),
				.b8(W2H22D),
				.c(c2D21H)
);

ninexnine_unit ninexnine_unit_5538(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2H00E),
				.b1(W2H01E),
				.b2(W2H02E),
				.b3(W2H10E),
				.b4(W2H11E),
				.b5(W2H12E),
				.b6(W2H20E),
				.b7(W2H21E),
				.b8(W2H22E),
				.c(c2E21H)
);

ninexnine_unit ninexnine_unit_5539(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2H00F),
				.b1(W2H01F),
				.b2(W2H02F),
				.b3(W2H10F),
				.b4(W2H11F),
				.b5(W2H12F),
				.b6(W2H20F),
				.b7(W2H21F),
				.b8(W2H22F),
				.c(c2F21H)
);

assign C221H=c2021H+c2121H+c2221H+c2321H+c2421H+c2521H+c2621H+c2721H+c2821H+c2921H+c2A21H+c2B21H+c2C21H+c2D21H+c2E21H+c2F21H;
assign A221H=(C221H>=0)?1:0;

assign P321H=A221H;

ninexnine_unit ninexnine_unit_5540(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2H000),
				.b1(W2H010),
				.b2(W2H020),
				.b3(W2H100),
				.b4(W2H110),
				.b5(W2H120),
				.b6(W2H200),
				.b7(W2H210),
				.b8(W2H220),
				.c(c2022H)
);

ninexnine_unit ninexnine_unit_5541(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2H001),
				.b1(W2H011),
				.b2(W2H021),
				.b3(W2H101),
				.b4(W2H111),
				.b5(W2H121),
				.b6(W2H201),
				.b7(W2H211),
				.b8(W2H221),
				.c(c2122H)
);

ninexnine_unit ninexnine_unit_5542(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2H002),
				.b1(W2H012),
				.b2(W2H022),
				.b3(W2H102),
				.b4(W2H112),
				.b5(W2H122),
				.b6(W2H202),
				.b7(W2H212),
				.b8(W2H222),
				.c(c2222H)
);

ninexnine_unit ninexnine_unit_5543(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2H003),
				.b1(W2H013),
				.b2(W2H023),
				.b3(W2H103),
				.b4(W2H113),
				.b5(W2H123),
				.b6(W2H203),
				.b7(W2H213),
				.b8(W2H223),
				.c(c2322H)
);

ninexnine_unit ninexnine_unit_5544(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2H004),
				.b1(W2H014),
				.b2(W2H024),
				.b3(W2H104),
				.b4(W2H114),
				.b5(W2H124),
				.b6(W2H204),
				.b7(W2H214),
				.b8(W2H224),
				.c(c2422H)
);

ninexnine_unit ninexnine_unit_5545(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2H005),
				.b1(W2H015),
				.b2(W2H025),
				.b3(W2H105),
				.b4(W2H115),
				.b5(W2H125),
				.b6(W2H205),
				.b7(W2H215),
				.b8(W2H225),
				.c(c2522H)
);

ninexnine_unit ninexnine_unit_5546(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2H006),
				.b1(W2H016),
				.b2(W2H026),
				.b3(W2H106),
				.b4(W2H116),
				.b5(W2H126),
				.b6(W2H206),
				.b7(W2H216),
				.b8(W2H226),
				.c(c2622H)
);

ninexnine_unit ninexnine_unit_5547(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2H007),
				.b1(W2H017),
				.b2(W2H027),
				.b3(W2H107),
				.b4(W2H117),
				.b5(W2H127),
				.b6(W2H207),
				.b7(W2H217),
				.b8(W2H227),
				.c(c2722H)
);

ninexnine_unit ninexnine_unit_5548(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2H008),
				.b1(W2H018),
				.b2(W2H028),
				.b3(W2H108),
				.b4(W2H118),
				.b5(W2H128),
				.b6(W2H208),
				.b7(W2H218),
				.b8(W2H228),
				.c(c2822H)
);

ninexnine_unit ninexnine_unit_5549(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2H009),
				.b1(W2H019),
				.b2(W2H029),
				.b3(W2H109),
				.b4(W2H119),
				.b5(W2H129),
				.b6(W2H209),
				.b7(W2H219),
				.b8(W2H229),
				.c(c2922H)
);

ninexnine_unit ninexnine_unit_5550(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2H00A),
				.b1(W2H01A),
				.b2(W2H02A),
				.b3(W2H10A),
				.b4(W2H11A),
				.b5(W2H12A),
				.b6(W2H20A),
				.b7(W2H21A),
				.b8(W2H22A),
				.c(c2A22H)
);

ninexnine_unit ninexnine_unit_5551(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2H00B),
				.b1(W2H01B),
				.b2(W2H02B),
				.b3(W2H10B),
				.b4(W2H11B),
				.b5(W2H12B),
				.b6(W2H20B),
				.b7(W2H21B),
				.b8(W2H22B),
				.c(c2B22H)
);

ninexnine_unit ninexnine_unit_5552(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2H00C),
				.b1(W2H01C),
				.b2(W2H02C),
				.b3(W2H10C),
				.b4(W2H11C),
				.b5(W2H12C),
				.b6(W2H20C),
				.b7(W2H21C),
				.b8(W2H22C),
				.c(c2C22H)
);

ninexnine_unit ninexnine_unit_5553(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2H00D),
				.b1(W2H01D),
				.b2(W2H02D),
				.b3(W2H10D),
				.b4(W2H11D),
				.b5(W2H12D),
				.b6(W2H20D),
				.b7(W2H21D),
				.b8(W2H22D),
				.c(c2D22H)
);

ninexnine_unit ninexnine_unit_5554(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2H00E),
				.b1(W2H01E),
				.b2(W2H02E),
				.b3(W2H10E),
				.b4(W2H11E),
				.b5(W2H12E),
				.b6(W2H20E),
				.b7(W2H21E),
				.b8(W2H22E),
				.c(c2E22H)
);

ninexnine_unit ninexnine_unit_5555(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2H00F),
				.b1(W2H01F),
				.b2(W2H02F),
				.b3(W2H10F),
				.b4(W2H11F),
				.b5(W2H12F),
				.b6(W2H20F),
				.b7(W2H21F),
				.b8(W2H22F),
				.c(c2F22H)
);

assign C222H=c2022H+c2122H+c2222H+c2322H+c2422H+c2522H+c2622H+c2722H+c2822H+c2922H+c2A22H+c2B22H+c2C22H+c2D22H+c2E22H+c2F22H;
assign A222H=(C222H>=0)?1:0;

assign P322H=A222H;

ninexnine_unit ninexnine_unit_5556(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2I000),
				.b1(W2I010),
				.b2(W2I020),
				.b3(W2I100),
				.b4(W2I110),
				.b5(W2I120),
				.b6(W2I200),
				.b7(W2I210),
				.b8(W2I220),
				.c(c2000I)
);

ninexnine_unit ninexnine_unit_5557(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2I001),
				.b1(W2I011),
				.b2(W2I021),
				.b3(W2I101),
				.b4(W2I111),
				.b5(W2I121),
				.b6(W2I201),
				.b7(W2I211),
				.b8(W2I221),
				.c(c2100I)
);

ninexnine_unit ninexnine_unit_5558(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2I002),
				.b1(W2I012),
				.b2(W2I022),
				.b3(W2I102),
				.b4(W2I112),
				.b5(W2I122),
				.b6(W2I202),
				.b7(W2I212),
				.b8(W2I222),
				.c(c2200I)
);

ninexnine_unit ninexnine_unit_5559(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2I003),
				.b1(W2I013),
				.b2(W2I023),
				.b3(W2I103),
				.b4(W2I113),
				.b5(W2I123),
				.b6(W2I203),
				.b7(W2I213),
				.b8(W2I223),
				.c(c2300I)
);

ninexnine_unit ninexnine_unit_5560(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2I004),
				.b1(W2I014),
				.b2(W2I024),
				.b3(W2I104),
				.b4(W2I114),
				.b5(W2I124),
				.b6(W2I204),
				.b7(W2I214),
				.b8(W2I224),
				.c(c2400I)
);

ninexnine_unit ninexnine_unit_5561(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2I005),
				.b1(W2I015),
				.b2(W2I025),
				.b3(W2I105),
				.b4(W2I115),
				.b5(W2I125),
				.b6(W2I205),
				.b7(W2I215),
				.b8(W2I225),
				.c(c2500I)
);

ninexnine_unit ninexnine_unit_5562(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2I006),
				.b1(W2I016),
				.b2(W2I026),
				.b3(W2I106),
				.b4(W2I116),
				.b5(W2I126),
				.b6(W2I206),
				.b7(W2I216),
				.b8(W2I226),
				.c(c2600I)
);

ninexnine_unit ninexnine_unit_5563(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2I007),
				.b1(W2I017),
				.b2(W2I027),
				.b3(W2I107),
				.b4(W2I117),
				.b5(W2I127),
				.b6(W2I207),
				.b7(W2I217),
				.b8(W2I227),
				.c(c2700I)
);

ninexnine_unit ninexnine_unit_5564(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2I008),
				.b1(W2I018),
				.b2(W2I028),
				.b3(W2I108),
				.b4(W2I118),
				.b5(W2I128),
				.b6(W2I208),
				.b7(W2I218),
				.b8(W2I228),
				.c(c2800I)
);

ninexnine_unit ninexnine_unit_5565(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2I009),
				.b1(W2I019),
				.b2(W2I029),
				.b3(W2I109),
				.b4(W2I119),
				.b5(W2I129),
				.b6(W2I209),
				.b7(W2I219),
				.b8(W2I229),
				.c(c2900I)
);

ninexnine_unit ninexnine_unit_5566(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2I00A),
				.b1(W2I01A),
				.b2(W2I02A),
				.b3(W2I10A),
				.b4(W2I11A),
				.b5(W2I12A),
				.b6(W2I20A),
				.b7(W2I21A),
				.b8(W2I22A),
				.c(c2A00I)
);

ninexnine_unit ninexnine_unit_5567(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2I00B),
				.b1(W2I01B),
				.b2(W2I02B),
				.b3(W2I10B),
				.b4(W2I11B),
				.b5(W2I12B),
				.b6(W2I20B),
				.b7(W2I21B),
				.b8(W2I22B),
				.c(c2B00I)
);

ninexnine_unit ninexnine_unit_5568(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2I00C),
				.b1(W2I01C),
				.b2(W2I02C),
				.b3(W2I10C),
				.b4(W2I11C),
				.b5(W2I12C),
				.b6(W2I20C),
				.b7(W2I21C),
				.b8(W2I22C),
				.c(c2C00I)
);

ninexnine_unit ninexnine_unit_5569(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2I00D),
				.b1(W2I01D),
				.b2(W2I02D),
				.b3(W2I10D),
				.b4(W2I11D),
				.b5(W2I12D),
				.b6(W2I20D),
				.b7(W2I21D),
				.b8(W2I22D),
				.c(c2D00I)
);

ninexnine_unit ninexnine_unit_5570(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2I00E),
				.b1(W2I01E),
				.b2(W2I02E),
				.b3(W2I10E),
				.b4(W2I11E),
				.b5(W2I12E),
				.b6(W2I20E),
				.b7(W2I21E),
				.b8(W2I22E),
				.c(c2E00I)
);

ninexnine_unit ninexnine_unit_5571(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2I00F),
				.b1(W2I01F),
				.b2(W2I02F),
				.b3(W2I10F),
				.b4(W2I11F),
				.b5(W2I12F),
				.b6(W2I20F),
				.b7(W2I21F),
				.b8(W2I22F),
				.c(c2F00I)
);

assign C200I=c2000I+c2100I+c2200I+c2300I+c2400I+c2500I+c2600I+c2700I+c2800I+c2900I+c2A00I+c2B00I+c2C00I+c2D00I+c2E00I+c2F00I;
assign A200I=(C200I>=0)?1:0;

assign P300I=A200I;

ninexnine_unit ninexnine_unit_5572(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2I000),
				.b1(W2I010),
				.b2(W2I020),
				.b3(W2I100),
				.b4(W2I110),
				.b5(W2I120),
				.b6(W2I200),
				.b7(W2I210),
				.b8(W2I220),
				.c(c2001I)
);

ninexnine_unit ninexnine_unit_5573(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2I001),
				.b1(W2I011),
				.b2(W2I021),
				.b3(W2I101),
				.b4(W2I111),
				.b5(W2I121),
				.b6(W2I201),
				.b7(W2I211),
				.b8(W2I221),
				.c(c2101I)
);

ninexnine_unit ninexnine_unit_5574(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2I002),
				.b1(W2I012),
				.b2(W2I022),
				.b3(W2I102),
				.b4(W2I112),
				.b5(W2I122),
				.b6(W2I202),
				.b7(W2I212),
				.b8(W2I222),
				.c(c2201I)
);

ninexnine_unit ninexnine_unit_5575(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2I003),
				.b1(W2I013),
				.b2(W2I023),
				.b3(W2I103),
				.b4(W2I113),
				.b5(W2I123),
				.b6(W2I203),
				.b7(W2I213),
				.b8(W2I223),
				.c(c2301I)
);

ninexnine_unit ninexnine_unit_5576(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2I004),
				.b1(W2I014),
				.b2(W2I024),
				.b3(W2I104),
				.b4(W2I114),
				.b5(W2I124),
				.b6(W2I204),
				.b7(W2I214),
				.b8(W2I224),
				.c(c2401I)
);

ninexnine_unit ninexnine_unit_5577(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2I005),
				.b1(W2I015),
				.b2(W2I025),
				.b3(W2I105),
				.b4(W2I115),
				.b5(W2I125),
				.b6(W2I205),
				.b7(W2I215),
				.b8(W2I225),
				.c(c2501I)
);

ninexnine_unit ninexnine_unit_5578(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2I006),
				.b1(W2I016),
				.b2(W2I026),
				.b3(W2I106),
				.b4(W2I116),
				.b5(W2I126),
				.b6(W2I206),
				.b7(W2I216),
				.b8(W2I226),
				.c(c2601I)
);

ninexnine_unit ninexnine_unit_5579(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2I007),
				.b1(W2I017),
				.b2(W2I027),
				.b3(W2I107),
				.b4(W2I117),
				.b5(W2I127),
				.b6(W2I207),
				.b7(W2I217),
				.b8(W2I227),
				.c(c2701I)
);

ninexnine_unit ninexnine_unit_5580(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2I008),
				.b1(W2I018),
				.b2(W2I028),
				.b3(W2I108),
				.b4(W2I118),
				.b5(W2I128),
				.b6(W2I208),
				.b7(W2I218),
				.b8(W2I228),
				.c(c2801I)
);

ninexnine_unit ninexnine_unit_5581(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2I009),
				.b1(W2I019),
				.b2(W2I029),
				.b3(W2I109),
				.b4(W2I119),
				.b5(W2I129),
				.b6(W2I209),
				.b7(W2I219),
				.b8(W2I229),
				.c(c2901I)
);

ninexnine_unit ninexnine_unit_5582(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2I00A),
				.b1(W2I01A),
				.b2(W2I02A),
				.b3(W2I10A),
				.b4(W2I11A),
				.b5(W2I12A),
				.b6(W2I20A),
				.b7(W2I21A),
				.b8(W2I22A),
				.c(c2A01I)
);

ninexnine_unit ninexnine_unit_5583(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2I00B),
				.b1(W2I01B),
				.b2(W2I02B),
				.b3(W2I10B),
				.b4(W2I11B),
				.b5(W2I12B),
				.b6(W2I20B),
				.b7(W2I21B),
				.b8(W2I22B),
				.c(c2B01I)
);

ninexnine_unit ninexnine_unit_5584(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2I00C),
				.b1(W2I01C),
				.b2(W2I02C),
				.b3(W2I10C),
				.b4(W2I11C),
				.b5(W2I12C),
				.b6(W2I20C),
				.b7(W2I21C),
				.b8(W2I22C),
				.c(c2C01I)
);

ninexnine_unit ninexnine_unit_5585(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2I00D),
				.b1(W2I01D),
				.b2(W2I02D),
				.b3(W2I10D),
				.b4(W2I11D),
				.b5(W2I12D),
				.b6(W2I20D),
				.b7(W2I21D),
				.b8(W2I22D),
				.c(c2D01I)
);

ninexnine_unit ninexnine_unit_5586(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2I00E),
				.b1(W2I01E),
				.b2(W2I02E),
				.b3(W2I10E),
				.b4(W2I11E),
				.b5(W2I12E),
				.b6(W2I20E),
				.b7(W2I21E),
				.b8(W2I22E),
				.c(c2E01I)
);

ninexnine_unit ninexnine_unit_5587(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2I00F),
				.b1(W2I01F),
				.b2(W2I02F),
				.b3(W2I10F),
				.b4(W2I11F),
				.b5(W2I12F),
				.b6(W2I20F),
				.b7(W2I21F),
				.b8(W2I22F),
				.c(c2F01I)
);

assign C201I=c2001I+c2101I+c2201I+c2301I+c2401I+c2501I+c2601I+c2701I+c2801I+c2901I+c2A01I+c2B01I+c2C01I+c2D01I+c2E01I+c2F01I;
assign A201I=(C201I>=0)?1:0;

assign P301I=A201I;

ninexnine_unit ninexnine_unit_5588(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2I000),
				.b1(W2I010),
				.b2(W2I020),
				.b3(W2I100),
				.b4(W2I110),
				.b5(W2I120),
				.b6(W2I200),
				.b7(W2I210),
				.b8(W2I220),
				.c(c2002I)
);

ninexnine_unit ninexnine_unit_5589(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2I001),
				.b1(W2I011),
				.b2(W2I021),
				.b3(W2I101),
				.b4(W2I111),
				.b5(W2I121),
				.b6(W2I201),
				.b7(W2I211),
				.b8(W2I221),
				.c(c2102I)
);

ninexnine_unit ninexnine_unit_5590(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2I002),
				.b1(W2I012),
				.b2(W2I022),
				.b3(W2I102),
				.b4(W2I112),
				.b5(W2I122),
				.b6(W2I202),
				.b7(W2I212),
				.b8(W2I222),
				.c(c2202I)
);

ninexnine_unit ninexnine_unit_5591(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2I003),
				.b1(W2I013),
				.b2(W2I023),
				.b3(W2I103),
				.b4(W2I113),
				.b5(W2I123),
				.b6(W2I203),
				.b7(W2I213),
				.b8(W2I223),
				.c(c2302I)
);

ninexnine_unit ninexnine_unit_5592(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2I004),
				.b1(W2I014),
				.b2(W2I024),
				.b3(W2I104),
				.b4(W2I114),
				.b5(W2I124),
				.b6(W2I204),
				.b7(W2I214),
				.b8(W2I224),
				.c(c2402I)
);

ninexnine_unit ninexnine_unit_5593(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2I005),
				.b1(W2I015),
				.b2(W2I025),
				.b3(W2I105),
				.b4(W2I115),
				.b5(W2I125),
				.b6(W2I205),
				.b7(W2I215),
				.b8(W2I225),
				.c(c2502I)
);

ninexnine_unit ninexnine_unit_5594(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2I006),
				.b1(W2I016),
				.b2(W2I026),
				.b3(W2I106),
				.b4(W2I116),
				.b5(W2I126),
				.b6(W2I206),
				.b7(W2I216),
				.b8(W2I226),
				.c(c2602I)
);

ninexnine_unit ninexnine_unit_5595(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2I007),
				.b1(W2I017),
				.b2(W2I027),
				.b3(W2I107),
				.b4(W2I117),
				.b5(W2I127),
				.b6(W2I207),
				.b7(W2I217),
				.b8(W2I227),
				.c(c2702I)
);

ninexnine_unit ninexnine_unit_5596(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2I008),
				.b1(W2I018),
				.b2(W2I028),
				.b3(W2I108),
				.b4(W2I118),
				.b5(W2I128),
				.b6(W2I208),
				.b7(W2I218),
				.b8(W2I228),
				.c(c2802I)
);

ninexnine_unit ninexnine_unit_5597(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2I009),
				.b1(W2I019),
				.b2(W2I029),
				.b3(W2I109),
				.b4(W2I119),
				.b5(W2I129),
				.b6(W2I209),
				.b7(W2I219),
				.b8(W2I229),
				.c(c2902I)
);

ninexnine_unit ninexnine_unit_5598(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2I00A),
				.b1(W2I01A),
				.b2(W2I02A),
				.b3(W2I10A),
				.b4(W2I11A),
				.b5(W2I12A),
				.b6(W2I20A),
				.b7(W2I21A),
				.b8(W2I22A),
				.c(c2A02I)
);

ninexnine_unit ninexnine_unit_5599(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2I00B),
				.b1(W2I01B),
				.b2(W2I02B),
				.b3(W2I10B),
				.b4(W2I11B),
				.b5(W2I12B),
				.b6(W2I20B),
				.b7(W2I21B),
				.b8(W2I22B),
				.c(c2B02I)
);

ninexnine_unit ninexnine_unit_5600(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2I00C),
				.b1(W2I01C),
				.b2(W2I02C),
				.b3(W2I10C),
				.b4(W2I11C),
				.b5(W2I12C),
				.b6(W2I20C),
				.b7(W2I21C),
				.b8(W2I22C),
				.c(c2C02I)
);

ninexnine_unit ninexnine_unit_5601(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2I00D),
				.b1(W2I01D),
				.b2(W2I02D),
				.b3(W2I10D),
				.b4(W2I11D),
				.b5(W2I12D),
				.b6(W2I20D),
				.b7(W2I21D),
				.b8(W2I22D),
				.c(c2D02I)
);

ninexnine_unit ninexnine_unit_5602(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2I00E),
				.b1(W2I01E),
				.b2(W2I02E),
				.b3(W2I10E),
				.b4(W2I11E),
				.b5(W2I12E),
				.b6(W2I20E),
				.b7(W2I21E),
				.b8(W2I22E),
				.c(c2E02I)
);

ninexnine_unit ninexnine_unit_5603(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2I00F),
				.b1(W2I01F),
				.b2(W2I02F),
				.b3(W2I10F),
				.b4(W2I11F),
				.b5(W2I12F),
				.b6(W2I20F),
				.b7(W2I21F),
				.b8(W2I22F),
				.c(c2F02I)
);

assign C202I=c2002I+c2102I+c2202I+c2302I+c2402I+c2502I+c2602I+c2702I+c2802I+c2902I+c2A02I+c2B02I+c2C02I+c2D02I+c2E02I+c2F02I;
assign A202I=(C202I>=0)?1:0;

assign P302I=A202I;

ninexnine_unit ninexnine_unit_5604(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2I000),
				.b1(W2I010),
				.b2(W2I020),
				.b3(W2I100),
				.b4(W2I110),
				.b5(W2I120),
				.b6(W2I200),
				.b7(W2I210),
				.b8(W2I220),
				.c(c2010I)
);

ninexnine_unit ninexnine_unit_5605(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2I001),
				.b1(W2I011),
				.b2(W2I021),
				.b3(W2I101),
				.b4(W2I111),
				.b5(W2I121),
				.b6(W2I201),
				.b7(W2I211),
				.b8(W2I221),
				.c(c2110I)
);

ninexnine_unit ninexnine_unit_5606(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2I002),
				.b1(W2I012),
				.b2(W2I022),
				.b3(W2I102),
				.b4(W2I112),
				.b5(W2I122),
				.b6(W2I202),
				.b7(W2I212),
				.b8(W2I222),
				.c(c2210I)
);

ninexnine_unit ninexnine_unit_5607(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2I003),
				.b1(W2I013),
				.b2(W2I023),
				.b3(W2I103),
				.b4(W2I113),
				.b5(W2I123),
				.b6(W2I203),
				.b7(W2I213),
				.b8(W2I223),
				.c(c2310I)
);

ninexnine_unit ninexnine_unit_5608(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2I004),
				.b1(W2I014),
				.b2(W2I024),
				.b3(W2I104),
				.b4(W2I114),
				.b5(W2I124),
				.b6(W2I204),
				.b7(W2I214),
				.b8(W2I224),
				.c(c2410I)
);

ninexnine_unit ninexnine_unit_5609(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2I005),
				.b1(W2I015),
				.b2(W2I025),
				.b3(W2I105),
				.b4(W2I115),
				.b5(W2I125),
				.b6(W2I205),
				.b7(W2I215),
				.b8(W2I225),
				.c(c2510I)
);

ninexnine_unit ninexnine_unit_5610(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2I006),
				.b1(W2I016),
				.b2(W2I026),
				.b3(W2I106),
				.b4(W2I116),
				.b5(W2I126),
				.b6(W2I206),
				.b7(W2I216),
				.b8(W2I226),
				.c(c2610I)
);

ninexnine_unit ninexnine_unit_5611(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2I007),
				.b1(W2I017),
				.b2(W2I027),
				.b3(W2I107),
				.b4(W2I117),
				.b5(W2I127),
				.b6(W2I207),
				.b7(W2I217),
				.b8(W2I227),
				.c(c2710I)
);

ninexnine_unit ninexnine_unit_5612(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2I008),
				.b1(W2I018),
				.b2(W2I028),
				.b3(W2I108),
				.b4(W2I118),
				.b5(W2I128),
				.b6(W2I208),
				.b7(W2I218),
				.b8(W2I228),
				.c(c2810I)
);

ninexnine_unit ninexnine_unit_5613(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2I009),
				.b1(W2I019),
				.b2(W2I029),
				.b3(W2I109),
				.b4(W2I119),
				.b5(W2I129),
				.b6(W2I209),
				.b7(W2I219),
				.b8(W2I229),
				.c(c2910I)
);

ninexnine_unit ninexnine_unit_5614(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2I00A),
				.b1(W2I01A),
				.b2(W2I02A),
				.b3(W2I10A),
				.b4(W2I11A),
				.b5(W2I12A),
				.b6(W2I20A),
				.b7(W2I21A),
				.b8(W2I22A),
				.c(c2A10I)
);

ninexnine_unit ninexnine_unit_5615(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2I00B),
				.b1(W2I01B),
				.b2(W2I02B),
				.b3(W2I10B),
				.b4(W2I11B),
				.b5(W2I12B),
				.b6(W2I20B),
				.b7(W2I21B),
				.b8(W2I22B),
				.c(c2B10I)
);

ninexnine_unit ninexnine_unit_5616(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2I00C),
				.b1(W2I01C),
				.b2(W2I02C),
				.b3(W2I10C),
				.b4(W2I11C),
				.b5(W2I12C),
				.b6(W2I20C),
				.b7(W2I21C),
				.b8(W2I22C),
				.c(c2C10I)
);

ninexnine_unit ninexnine_unit_5617(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2I00D),
				.b1(W2I01D),
				.b2(W2I02D),
				.b3(W2I10D),
				.b4(W2I11D),
				.b5(W2I12D),
				.b6(W2I20D),
				.b7(W2I21D),
				.b8(W2I22D),
				.c(c2D10I)
);

ninexnine_unit ninexnine_unit_5618(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2I00E),
				.b1(W2I01E),
				.b2(W2I02E),
				.b3(W2I10E),
				.b4(W2I11E),
				.b5(W2I12E),
				.b6(W2I20E),
				.b7(W2I21E),
				.b8(W2I22E),
				.c(c2E10I)
);

ninexnine_unit ninexnine_unit_5619(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2I00F),
				.b1(W2I01F),
				.b2(W2I02F),
				.b3(W2I10F),
				.b4(W2I11F),
				.b5(W2I12F),
				.b6(W2I20F),
				.b7(W2I21F),
				.b8(W2I22F),
				.c(c2F10I)
);

assign C210I=c2010I+c2110I+c2210I+c2310I+c2410I+c2510I+c2610I+c2710I+c2810I+c2910I+c2A10I+c2B10I+c2C10I+c2D10I+c2E10I+c2F10I;
assign A210I=(C210I>=0)?1:0;

assign P310I=A210I;

ninexnine_unit ninexnine_unit_5620(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2I000),
				.b1(W2I010),
				.b2(W2I020),
				.b3(W2I100),
				.b4(W2I110),
				.b5(W2I120),
				.b6(W2I200),
				.b7(W2I210),
				.b8(W2I220),
				.c(c2011I)
);

ninexnine_unit ninexnine_unit_5621(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2I001),
				.b1(W2I011),
				.b2(W2I021),
				.b3(W2I101),
				.b4(W2I111),
				.b5(W2I121),
				.b6(W2I201),
				.b7(W2I211),
				.b8(W2I221),
				.c(c2111I)
);

ninexnine_unit ninexnine_unit_5622(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2I002),
				.b1(W2I012),
				.b2(W2I022),
				.b3(W2I102),
				.b4(W2I112),
				.b5(W2I122),
				.b6(W2I202),
				.b7(W2I212),
				.b8(W2I222),
				.c(c2211I)
);

ninexnine_unit ninexnine_unit_5623(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2I003),
				.b1(W2I013),
				.b2(W2I023),
				.b3(W2I103),
				.b4(W2I113),
				.b5(W2I123),
				.b6(W2I203),
				.b7(W2I213),
				.b8(W2I223),
				.c(c2311I)
);

ninexnine_unit ninexnine_unit_5624(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2I004),
				.b1(W2I014),
				.b2(W2I024),
				.b3(W2I104),
				.b4(W2I114),
				.b5(W2I124),
				.b6(W2I204),
				.b7(W2I214),
				.b8(W2I224),
				.c(c2411I)
);

ninexnine_unit ninexnine_unit_5625(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2I005),
				.b1(W2I015),
				.b2(W2I025),
				.b3(W2I105),
				.b4(W2I115),
				.b5(W2I125),
				.b6(W2I205),
				.b7(W2I215),
				.b8(W2I225),
				.c(c2511I)
);

ninexnine_unit ninexnine_unit_5626(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2I006),
				.b1(W2I016),
				.b2(W2I026),
				.b3(W2I106),
				.b4(W2I116),
				.b5(W2I126),
				.b6(W2I206),
				.b7(W2I216),
				.b8(W2I226),
				.c(c2611I)
);

ninexnine_unit ninexnine_unit_5627(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2I007),
				.b1(W2I017),
				.b2(W2I027),
				.b3(W2I107),
				.b4(W2I117),
				.b5(W2I127),
				.b6(W2I207),
				.b7(W2I217),
				.b8(W2I227),
				.c(c2711I)
);

ninexnine_unit ninexnine_unit_5628(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2I008),
				.b1(W2I018),
				.b2(W2I028),
				.b3(W2I108),
				.b4(W2I118),
				.b5(W2I128),
				.b6(W2I208),
				.b7(W2I218),
				.b8(W2I228),
				.c(c2811I)
);

ninexnine_unit ninexnine_unit_5629(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2I009),
				.b1(W2I019),
				.b2(W2I029),
				.b3(W2I109),
				.b4(W2I119),
				.b5(W2I129),
				.b6(W2I209),
				.b7(W2I219),
				.b8(W2I229),
				.c(c2911I)
);

ninexnine_unit ninexnine_unit_5630(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2I00A),
				.b1(W2I01A),
				.b2(W2I02A),
				.b3(W2I10A),
				.b4(W2I11A),
				.b5(W2I12A),
				.b6(W2I20A),
				.b7(W2I21A),
				.b8(W2I22A),
				.c(c2A11I)
);

ninexnine_unit ninexnine_unit_5631(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2I00B),
				.b1(W2I01B),
				.b2(W2I02B),
				.b3(W2I10B),
				.b4(W2I11B),
				.b5(W2I12B),
				.b6(W2I20B),
				.b7(W2I21B),
				.b8(W2I22B),
				.c(c2B11I)
);

ninexnine_unit ninexnine_unit_5632(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2I00C),
				.b1(W2I01C),
				.b2(W2I02C),
				.b3(W2I10C),
				.b4(W2I11C),
				.b5(W2I12C),
				.b6(W2I20C),
				.b7(W2I21C),
				.b8(W2I22C),
				.c(c2C11I)
);

ninexnine_unit ninexnine_unit_5633(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2I00D),
				.b1(W2I01D),
				.b2(W2I02D),
				.b3(W2I10D),
				.b4(W2I11D),
				.b5(W2I12D),
				.b6(W2I20D),
				.b7(W2I21D),
				.b8(W2I22D),
				.c(c2D11I)
);

ninexnine_unit ninexnine_unit_5634(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2I00E),
				.b1(W2I01E),
				.b2(W2I02E),
				.b3(W2I10E),
				.b4(W2I11E),
				.b5(W2I12E),
				.b6(W2I20E),
				.b7(W2I21E),
				.b8(W2I22E),
				.c(c2E11I)
);

ninexnine_unit ninexnine_unit_5635(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2I00F),
				.b1(W2I01F),
				.b2(W2I02F),
				.b3(W2I10F),
				.b4(W2I11F),
				.b5(W2I12F),
				.b6(W2I20F),
				.b7(W2I21F),
				.b8(W2I22F),
				.c(c2F11I)
);

assign C211I=c2011I+c2111I+c2211I+c2311I+c2411I+c2511I+c2611I+c2711I+c2811I+c2911I+c2A11I+c2B11I+c2C11I+c2D11I+c2E11I+c2F11I;
assign A211I=(C211I>=0)?1:0;

assign P311I=A211I;

ninexnine_unit ninexnine_unit_5636(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2I000),
				.b1(W2I010),
				.b2(W2I020),
				.b3(W2I100),
				.b4(W2I110),
				.b5(W2I120),
				.b6(W2I200),
				.b7(W2I210),
				.b8(W2I220),
				.c(c2012I)
);

ninexnine_unit ninexnine_unit_5637(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2I001),
				.b1(W2I011),
				.b2(W2I021),
				.b3(W2I101),
				.b4(W2I111),
				.b5(W2I121),
				.b6(W2I201),
				.b7(W2I211),
				.b8(W2I221),
				.c(c2112I)
);

ninexnine_unit ninexnine_unit_5638(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2I002),
				.b1(W2I012),
				.b2(W2I022),
				.b3(W2I102),
				.b4(W2I112),
				.b5(W2I122),
				.b6(W2I202),
				.b7(W2I212),
				.b8(W2I222),
				.c(c2212I)
);

ninexnine_unit ninexnine_unit_5639(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2I003),
				.b1(W2I013),
				.b2(W2I023),
				.b3(W2I103),
				.b4(W2I113),
				.b5(W2I123),
				.b6(W2I203),
				.b7(W2I213),
				.b8(W2I223),
				.c(c2312I)
);

ninexnine_unit ninexnine_unit_5640(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2I004),
				.b1(W2I014),
				.b2(W2I024),
				.b3(W2I104),
				.b4(W2I114),
				.b5(W2I124),
				.b6(W2I204),
				.b7(W2I214),
				.b8(W2I224),
				.c(c2412I)
);

ninexnine_unit ninexnine_unit_5641(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2I005),
				.b1(W2I015),
				.b2(W2I025),
				.b3(W2I105),
				.b4(W2I115),
				.b5(W2I125),
				.b6(W2I205),
				.b7(W2I215),
				.b8(W2I225),
				.c(c2512I)
);

ninexnine_unit ninexnine_unit_5642(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2I006),
				.b1(W2I016),
				.b2(W2I026),
				.b3(W2I106),
				.b4(W2I116),
				.b5(W2I126),
				.b6(W2I206),
				.b7(W2I216),
				.b8(W2I226),
				.c(c2612I)
);

ninexnine_unit ninexnine_unit_5643(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2I007),
				.b1(W2I017),
				.b2(W2I027),
				.b3(W2I107),
				.b4(W2I117),
				.b5(W2I127),
				.b6(W2I207),
				.b7(W2I217),
				.b8(W2I227),
				.c(c2712I)
);

ninexnine_unit ninexnine_unit_5644(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2I008),
				.b1(W2I018),
				.b2(W2I028),
				.b3(W2I108),
				.b4(W2I118),
				.b5(W2I128),
				.b6(W2I208),
				.b7(W2I218),
				.b8(W2I228),
				.c(c2812I)
);

ninexnine_unit ninexnine_unit_5645(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2I009),
				.b1(W2I019),
				.b2(W2I029),
				.b3(W2I109),
				.b4(W2I119),
				.b5(W2I129),
				.b6(W2I209),
				.b7(W2I219),
				.b8(W2I229),
				.c(c2912I)
);

ninexnine_unit ninexnine_unit_5646(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2I00A),
				.b1(W2I01A),
				.b2(W2I02A),
				.b3(W2I10A),
				.b4(W2I11A),
				.b5(W2I12A),
				.b6(W2I20A),
				.b7(W2I21A),
				.b8(W2I22A),
				.c(c2A12I)
);

ninexnine_unit ninexnine_unit_5647(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2I00B),
				.b1(W2I01B),
				.b2(W2I02B),
				.b3(W2I10B),
				.b4(W2I11B),
				.b5(W2I12B),
				.b6(W2I20B),
				.b7(W2I21B),
				.b8(W2I22B),
				.c(c2B12I)
);

ninexnine_unit ninexnine_unit_5648(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2I00C),
				.b1(W2I01C),
				.b2(W2I02C),
				.b3(W2I10C),
				.b4(W2I11C),
				.b5(W2I12C),
				.b6(W2I20C),
				.b7(W2I21C),
				.b8(W2I22C),
				.c(c2C12I)
);

ninexnine_unit ninexnine_unit_5649(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2I00D),
				.b1(W2I01D),
				.b2(W2I02D),
				.b3(W2I10D),
				.b4(W2I11D),
				.b5(W2I12D),
				.b6(W2I20D),
				.b7(W2I21D),
				.b8(W2I22D),
				.c(c2D12I)
);

ninexnine_unit ninexnine_unit_5650(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2I00E),
				.b1(W2I01E),
				.b2(W2I02E),
				.b3(W2I10E),
				.b4(W2I11E),
				.b5(W2I12E),
				.b6(W2I20E),
				.b7(W2I21E),
				.b8(W2I22E),
				.c(c2E12I)
);

ninexnine_unit ninexnine_unit_5651(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2I00F),
				.b1(W2I01F),
				.b2(W2I02F),
				.b3(W2I10F),
				.b4(W2I11F),
				.b5(W2I12F),
				.b6(W2I20F),
				.b7(W2I21F),
				.b8(W2I22F),
				.c(c2F12I)
);

assign C212I=c2012I+c2112I+c2212I+c2312I+c2412I+c2512I+c2612I+c2712I+c2812I+c2912I+c2A12I+c2B12I+c2C12I+c2D12I+c2E12I+c2F12I;
assign A212I=(C212I>=0)?1:0;

assign P312I=A212I;

ninexnine_unit ninexnine_unit_5652(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2I000),
				.b1(W2I010),
				.b2(W2I020),
				.b3(W2I100),
				.b4(W2I110),
				.b5(W2I120),
				.b6(W2I200),
				.b7(W2I210),
				.b8(W2I220),
				.c(c2020I)
);

ninexnine_unit ninexnine_unit_5653(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2I001),
				.b1(W2I011),
				.b2(W2I021),
				.b3(W2I101),
				.b4(W2I111),
				.b5(W2I121),
				.b6(W2I201),
				.b7(W2I211),
				.b8(W2I221),
				.c(c2120I)
);

ninexnine_unit ninexnine_unit_5654(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2I002),
				.b1(W2I012),
				.b2(W2I022),
				.b3(W2I102),
				.b4(W2I112),
				.b5(W2I122),
				.b6(W2I202),
				.b7(W2I212),
				.b8(W2I222),
				.c(c2220I)
);

ninexnine_unit ninexnine_unit_5655(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2I003),
				.b1(W2I013),
				.b2(W2I023),
				.b3(W2I103),
				.b4(W2I113),
				.b5(W2I123),
				.b6(W2I203),
				.b7(W2I213),
				.b8(W2I223),
				.c(c2320I)
);

ninexnine_unit ninexnine_unit_5656(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2I004),
				.b1(W2I014),
				.b2(W2I024),
				.b3(W2I104),
				.b4(W2I114),
				.b5(W2I124),
				.b6(W2I204),
				.b7(W2I214),
				.b8(W2I224),
				.c(c2420I)
);

ninexnine_unit ninexnine_unit_5657(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2I005),
				.b1(W2I015),
				.b2(W2I025),
				.b3(W2I105),
				.b4(W2I115),
				.b5(W2I125),
				.b6(W2I205),
				.b7(W2I215),
				.b8(W2I225),
				.c(c2520I)
);

ninexnine_unit ninexnine_unit_5658(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2I006),
				.b1(W2I016),
				.b2(W2I026),
				.b3(W2I106),
				.b4(W2I116),
				.b5(W2I126),
				.b6(W2I206),
				.b7(W2I216),
				.b8(W2I226),
				.c(c2620I)
);

ninexnine_unit ninexnine_unit_5659(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2I007),
				.b1(W2I017),
				.b2(W2I027),
				.b3(W2I107),
				.b4(W2I117),
				.b5(W2I127),
				.b6(W2I207),
				.b7(W2I217),
				.b8(W2I227),
				.c(c2720I)
);

ninexnine_unit ninexnine_unit_5660(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2I008),
				.b1(W2I018),
				.b2(W2I028),
				.b3(W2I108),
				.b4(W2I118),
				.b5(W2I128),
				.b6(W2I208),
				.b7(W2I218),
				.b8(W2I228),
				.c(c2820I)
);

ninexnine_unit ninexnine_unit_5661(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2I009),
				.b1(W2I019),
				.b2(W2I029),
				.b3(W2I109),
				.b4(W2I119),
				.b5(W2I129),
				.b6(W2I209),
				.b7(W2I219),
				.b8(W2I229),
				.c(c2920I)
);

ninexnine_unit ninexnine_unit_5662(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2I00A),
				.b1(W2I01A),
				.b2(W2I02A),
				.b3(W2I10A),
				.b4(W2I11A),
				.b5(W2I12A),
				.b6(W2I20A),
				.b7(W2I21A),
				.b8(W2I22A),
				.c(c2A20I)
);

ninexnine_unit ninexnine_unit_5663(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2I00B),
				.b1(W2I01B),
				.b2(W2I02B),
				.b3(W2I10B),
				.b4(W2I11B),
				.b5(W2I12B),
				.b6(W2I20B),
				.b7(W2I21B),
				.b8(W2I22B),
				.c(c2B20I)
);

ninexnine_unit ninexnine_unit_5664(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2I00C),
				.b1(W2I01C),
				.b2(W2I02C),
				.b3(W2I10C),
				.b4(W2I11C),
				.b5(W2I12C),
				.b6(W2I20C),
				.b7(W2I21C),
				.b8(W2I22C),
				.c(c2C20I)
);

ninexnine_unit ninexnine_unit_5665(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2I00D),
				.b1(W2I01D),
				.b2(W2I02D),
				.b3(W2I10D),
				.b4(W2I11D),
				.b5(W2I12D),
				.b6(W2I20D),
				.b7(W2I21D),
				.b8(W2I22D),
				.c(c2D20I)
);

ninexnine_unit ninexnine_unit_5666(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2I00E),
				.b1(W2I01E),
				.b2(W2I02E),
				.b3(W2I10E),
				.b4(W2I11E),
				.b5(W2I12E),
				.b6(W2I20E),
				.b7(W2I21E),
				.b8(W2I22E),
				.c(c2E20I)
);

ninexnine_unit ninexnine_unit_5667(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2I00F),
				.b1(W2I01F),
				.b2(W2I02F),
				.b3(W2I10F),
				.b4(W2I11F),
				.b5(W2I12F),
				.b6(W2I20F),
				.b7(W2I21F),
				.b8(W2I22F),
				.c(c2F20I)
);

assign C220I=c2020I+c2120I+c2220I+c2320I+c2420I+c2520I+c2620I+c2720I+c2820I+c2920I+c2A20I+c2B20I+c2C20I+c2D20I+c2E20I+c2F20I;
assign A220I=(C220I>=0)?1:0;

assign P320I=A220I;

ninexnine_unit ninexnine_unit_5668(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2I000),
				.b1(W2I010),
				.b2(W2I020),
				.b3(W2I100),
				.b4(W2I110),
				.b5(W2I120),
				.b6(W2I200),
				.b7(W2I210),
				.b8(W2I220),
				.c(c2021I)
);

ninexnine_unit ninexnine_unit_5669(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2I001),
				.b1(W2I011),
				.b2(W2I021),
				.b3(W2I101),
				.b4(W2I111),
				.b5(W2I121),
				.b6(W2I201),
				.b7(W2I211),
				.b8(W2I221),
				.c(c2121I)
);

ninexnine_unit ninexnine_unit_5670(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2I002),
				.b1(W2I012),
				.b2(W2I022),
				.b3(W2I102),
				.b4(W2I112),
				.b5(W2I122),
				.b6(W2I202),
				.b7(W2I212),
				.b8(W2I222),
				.c(c2221I)
);

ninexnine_unit ninexnine_unit_5671(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2I003),
				.b1(W2I013),
				.b2(W2I023),
				.b3(W2I103),
				.b4(W2I113),
				.b5(W2I123),
				.b6(W2I203),
				.b7(W2I213),
				.b8(W2I223),
				.c(c2321I)
);

ninexnine_unit ninexnine_unit_5672(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2I004),
				.b1(W2I014),
				.b2(W2I024),
				.b3(W2I104),
				.b4(W2I114),
				.b5(W2I124),
				.b6(W2I204),
				.b7(W2I214),
				.b8(W2I224),
				.c(c2421I)
);

ninexnine_unit ninexnine_unit_5673(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2I005),
				.b1(W2I015),
				.b2(W2I025),
				.b3(W2I105),
				.b4(W2I115),
				.b5(W2I125),
				.b6(W2I205),
				.b7(W2I215),
				.b8(W2I225),
				.c(c2521I)
);

ninexnine_unit ninexnine_unit_5674(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2I006),
				.b1(W2I016),
				.b2(W2I026),
				.b3(W2I106),
				.b4(W2I116),
				.b5(W2I126),
				.b6(W2I206),
				.b7(W2I216),
				.b8(W2I226),
				.c(c2621I)
);

ninexnine_unit ninexnine_unit_5675(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2I007),
				.b1(W2I017),
				.b2(W2I027),
				.b3(W2I107),
				.b4(W2I117),
				.b5(W2I127),
				.b6(W2I207),
				.b7(W2I217),
				.b8(W2I227),
				.c(c2721I)
);

ninexnine_unit ninexnine_unit_5676(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2I008),
				.b1(W2I018),
				.b2(W2I028),
				.b3(W2I108),
				.b4(W2I118),
				.b5(W2I128),
				.b6(W2I208),
				.b7(W2I218),
				.b8(W2I228),
				.c(c2821I)
);

ninexnine_unit ninexnine_unit_5677(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2I009),
				.b1(W2I019),
				.b2(W2I029),
				.b3(W2I109),
				.b4(W2I119),
				.b5(W2I129),
				.b6(W2I209),
				.b7(W2I219),
				.b8(W2I229),
				.c(c2921I)
);

ninexnine_unit ninexnine_unit_5678(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2I00A),
				.b1(W2I01A),
				.b2(W2I02A),
				.b3(W2I10A),
				.b4(W2I11A),
				.b5(W2I12A),
				.b6(W2I20A),
				.b7(W2I21A),
				.b8(W2I22A),
				.c(c2A21I)
);

ninexnine_unit ninexnine_unit_5679(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2I00B),
				.b1(W2I01B),
				.b2(W2I02B),
				.b3(W2I10B),
				.b4(W2I11B),
				.b5(W2I12B),
				.b6(W2I20B),
				.b7(W2I21B),
				.b8(W2I22B),
				.c(c2B21I)
);

ninexnine_unit ninexnine_unit_5680(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2I00C),
				.b1(W2I01C),
				.b2(W2I02C),
				.b3(W2I10C),
				.b4(W2I11C),
				.b5(W2I12C),
				.b6(W2I20C),
				.b7(W2I21C),
				.b8(W2I22C),
				.c(c2C21I)
);

ninexnine_unit ninexnine_unit_5681(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2I00D),
				.b1(W2I01D),
				.b2(W2I02D),
				.b3(W2I10D),
				.b4(W2I11D),
				.b5(W2I12D),
				.b6(W2I20D),
				.b7(W2I21D),
				.b8(W2I22D),
				.c(c2D21I)
);

ninexnine_unit ninexnine_unit_5682(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2I00E),
				.b1(W2I01E),
				.b2(W2I02E),
				.b3(W2I10E),
				.b4(W2I11E),
				.b5(W2I12E),
				.b6(W2I20E),
				.b7(W2I21E),
				.b8(W2I22E),
				.c(c2E21I)
);

ninexnine_unit ninexnine_unit_5683(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2I00F),
				.b1(W2I01F),
				.b2(W2I02F),
				.b3(W2I10F),
				.b4(W2I11F),
				.b5(W2I12F),
				.b6(W2I20F),
				.b7(W2I21F),
				.b8(W2I22F),
				.c(c2F21I)
);

assign C221I=c2021I+c2121I+c2221I+c2321I+c2421I+c2521I+c2621I+c2721I+c2821I+c2921I+c2A21I+c2B21I+c2C21I+c2D21I+c2E21I+c2F21I;
assign A221I=(C221I>=0)?1:0;

assign P321I=A221I;

ninexnine_unit ninexnine_unit_5684(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2I000),
				.b1(W2I010),
				.b2(W2I020),
				.b3(W2I100),
				.b4(W2I110),
				.b5(W2I120),
				.b6(W2I200),
				.b7(W2I210),
				.b8(W2I220),
				.c(c2022I)
);

ninexnine_unit ninexnine_unit_5685(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2I001),
				.b1(W2I011),
				.b2(W2I021),
				.b3(W2I101),
				.b4(W2I111),
				.b5(W2I121),
				.b6(W2I201),
				.b7(W2I211),
				.b8(W2I221),
				.c(c2122I)
);

ninexnine_unit ninexnine_unit_5686(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2I002),
				.b1(W2I012),
				.b2(W2I022),
				.b3(W2I102),
				.b4(W2I112),
				.b5(W2I122),
				.b6(W2I202),
				.b7(W2I212),
				.b8(W2I222),
				.c(c2222I)
);

ninexnine_unit ninexnine_unit_5687(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2I003),
				.b1(W2I013),
				.b2(W2I023),
				.b3(W2I103),
				.b4(W2I113),
				.b5(W2I123),
				.b6(W2I203),
				.b7(W2I213),
				.b8(W2I223),
				.c(c2322I)
);

ninexnine_unit ninexnine_unit_5688(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2I004),
				.b1(W2I014),
				.b2(W2I024),
				.b3(W2I104),
				.b4(W2I114),
				.b5(W2I124),
				.b6(W2I204),
				.b7(W2I214),
				.b8(W2I224),
				.c(c2422I)
);

ninexnine_unit ninexnine_unit_5689(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2I005),
				.b1(W2I015),
				.b2(W2I025),
				.b3(W2I105),
				.b4(W2I115),
				.b5(W2I125),
				.b6(W2I205),
				.b7(W2I215),
				.b8(W2I225),
				.c(c2522I)
);

ninexnine_unit ninexnine_unit_5690(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2I006),
				.b1(W2I016),
				.b2(W2I026),
				.b3(W2I106),
				.b4(W2I116),
				.b5(W2I126),
				.b6(W2I206),
				.b7(W2I216),
				.b8(W2I226),
				.c(c2622I)
);

ninexnine_unit ninexnine_unit_5691(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2I007),
				.b1(W2I017),
				.b2(W2I027),
				.b3(W2I107),
				.b4(W2I117),
				.b5(W2I127),
				.b6(W2I207),
				.b7(W2I217),
				.b8(W2I227),
				.c(c2722I)
);

ninexnine_unit ninexnine_unit_5692(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2I008),
				.b1(W2I018),
				.b2(W2I028),
				.b3(W2I108),
				.b4(W2I118),
				.b5(W2I128),
				.b6(W2I208),
				.b7(W2I218),
				.b8(W2I228),
				.c(c2822I)
);

ninexnine_unit ninexnine_unit_5693(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2I009),
				.b1(W2I019),
				.b2(W2I029),
				.b3(W2I109),
				.b4(W2I119),
				.b5(W2I129),
				.b6(W2I209),
				.b7(W2I219),
				.b8(W2I229),
				.c(c2922I)
);

ninexnine_unit ninexnine_unit_5694(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2I00A),
				.b1(W2I01A),
				.b2(W2I02A),
				.b3(W2I10A),
				.b4(W2I11A),
				.b5(W2I12A),
				.b6(W2I20A),
				.b7(W2I21A),
				.b8(W2I22A),
				.c(c2A22I)
);

ninexnine_unit ninexnine_unit_5695(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2I00B),
				.b1(W2I01B),
				.b2(W2I02B),
				.b3(W2I10B),
				.b4(W2I11B),
				.b5(W2I12B),
				.b6(W2I20B),
				.b7(W2I21B),
				.b8(W2I22B),
				.c(c2B22I)
);

ninexnine_unit ninexnine_unit_5696(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2I00C),
				.b1(W2I01C),
				.b2(W2I02C),
				.b3(W2I10C),
				.b4(W2I11C),
				.b5(W2I12C),
				.b6(W2I20C),
				.b7(W2I21C),
				.b8(W2I22C),
				.c(c2C22I)
);

ninexnine_unit ninexnine_unit_5697(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2I00D),
				.b1(W2I01D),
				.b2(W2I02D),
				.b3(W2I10D),
				.b4(W2I11D),
				.b5(W2I12D),
				.b6(W2I20D),
				.b7(W2I21D),
				.b8(W2I22D),
				.c(c2D22I)
);

ninexnine_unit ninexnine_unit_5698(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2I00E),
				.b1(W2I01E),
				.b2(W2I02E),
				.b3(W2I10E),
				.b4(W2I11E),
				.b5(W2I12E),
				.b6(W2I20E),
				.b7(W2I21E),
				.b8(W2I22E),
				.c(c2E22I)
);

ninexnine_unit ninexnine_unit_5699(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2I00F),
				.b1(W2I01F),
				.b2(W2I02F),
				.b3(W2I10F),
				.b4(W2I11F),
				.b5(W2I12F),
				.b6(W2I20F),
				.b7(W2I21F),
				.b8(W2I22F),
				.c(c2F22I)
);

assign C222I=c2022I+c2122I+c2222I+c2322I+c2422I+c2522I+c2622I+c2722I+c2822I+c2922I+c2A22I+c2B22I+c2C22I+c2D22I+c2E22I+c2F22I;
assign A222I=(C222I>=0)?1:0;

assign P322I=A222I;

ninexnine_unit ninexnine_unit_5700(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2J000),
				.b1(W2J010),
				.b2(W2J020),
				.b3(W2J100),
				.b4(W2J110),
				.b5(W2J120),
				.b6(W2J200),
				.b7(W2J210),
				.b8(W2J220),
				.c(c2000J)
);

ninexnine_unit ninexnine_unit_5701(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2J001),
				.b1(W2J011),
				.b2(W2J021),
				.b3(W2J101),
				.b4(W2J111),
				.b5(W2J121),
				.b6(W2J201),
				.b7(W2J211),
				.b8(W2J221),
				.c(c2100J)
);

ninexnine_unit ninexnine_unit_5702(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2J002),
				.b1(W2J012),
				.b2(W2J022),
				.b3(W2J102),
				.b4(W2J112),
				.b5(W2J122),
				.b6(W2J202),
				.b7(W2J212),
				.b8(W2J222),
				.c(c2200J)
);

ninexnine_unit ninexnine_unit_5703(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2J003),
				.b1(W2J013),
				.b2(W2J023),
				.b3(W2J103),
				.b4(W2J113),
				.b5(W2J123),
				.b6(W2J203),
				.b7(W2J213),
				.b8(W2J223),
				.c(c2300J)
);

ninexnine_unit ninexnine_unit_5704(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2J004),
				.b1(W2J014),
				.b2(W2J024),
				.b3(W2J104),
				.b4(W2J114),
				.b5(W2J124),
				.b6(W2J204),
				.b7(W2J214),
				.b8(W2J224),
				.c(c2400J)
);

ninexnine_unit ninexnine_unit_5705(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2J005),
				.b1(W2J015),
				.b2(W2J025),
				.b3(W2J105),
				.b4(W2J115),
				.b5(W2J125),
				.b6(W2J205),
				.b7(W2J215),
				.b8(W2J225),
				.c(c2500J)
);

ninexnine_unit ninexnine_unit_5706(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2J006),
				.b1(W2J016),
				.b2(W2J026),
				.b3(W2J106),
				.b4(W2J116),
				.b5(W2J126),
				.b6(W2J206),
				.b7(W2J216),
				.b8(W2J226),
				.c(c2600J)
);

ninexnine_unit ninexnine_unit_5707(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2J007),
				.b1(W2J017),
				.b2(W2J027),
				.b3(W2J107),
				.b4(W2J117),
				.b5(W2J127),
				.b6(W2J207),
				.b7(W2J217),
				.b8(W2J227),
				.c(c2700J)
);

ninexnine_unit ninexnine_unit_5708(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2J008),
				.b1(W2J018),
				.b2(W2J028),
				.b3(W2J108),
				.b4(W2J118),
				.b5(W2J128),
				.b6(W2J208),
				.b7(W2J218),
				.b8(W2J228),
				.c(c2800J)
);

ninexnine_unit ninexnine_unit_5709(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2J009),
				.b1(W2J019),
				.b2(W2J029),
				.b3(W2J109),
				.b4(W2J119),
				.b5(W2J129),
				.b6(W2J209),
				.b7(W2J219),
				.b8(W2J229),
				.c(c2900J)
);

ninexnine_unit ninexnine_unit_5710(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2J00A),
				.b1(W2J01A),
				.b2(W2J02A),
				.b3(W2J10A),
				.b4(W2J11A),
				.b5(W2J12A),
				.b6(W2J20A),
				.b7(W2J21A),
				.b8(W2J22A),
				.c(c2A00J)
);

ninexnine_unit ninexnine_unit_5711(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2J00B),
				.b1(W2J01B),
				.b2(W2J02B),
				.b3(W2J10B),
				.b4(W2J11B),
				.b5(W2J12B),
				.b6(W2J20B),
				.b7(W2J21B),
				.b8(W2J22B),
				.c(c2B00J)
);

ninexnine_unit ninexnine_unit_5712(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2J00C),
				.b1(W2J01C),
				.b2(W2J02C),
				.b3(W2J10C),
				.b4(W2J11C),
				.b5(W2J12C),
				.b6(W2J20C),
				.b7(W2J21C),
				.b8(W2J22C),
				.c(c2C00J)
);

ninexnine_unit ninexnine_unit_5713(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2J00D),
				.b1(W2J01D),
				.b2(W2J02D),
				.b3(W2J10D),
				.b4(W2J11D),
				.b5(W2J12D),
				.b6(W2J20D),
				.b7(W2J21D),
				.b8(W2J22D),
				.c(c2D00J)
);

ninexnine_unit ninexnine_unit_5714(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2J00E),
				.b1(W2J01E),
				.b2(W2J02E),
				.b3(W2J10E),
				.b4(W2J11E),
				.b5(W2J12E),
				.b6(W2J20E),
				.b7(W2J21E),
				.b8(W2J22E),
				.c(c2E00J)
);

ninexnine_unit ninexnine_unit_5715(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2J00F),
				.b1(W2J01F),
				.b2(W2J02F),
				.b3(W2J10F),
				.b4(W2J11F),
				.b5(W2J12F),
				.b6(W2J20F),
				.b7(W2J21F),
				.b8(W2J22F),
				.c(c2F00J)
);

assign C200J=c2000J+c2100J+c2200J+c2300J+c2400J+c2500J+c2600J+c2700J+c2800J+c2900J+c2A00J+c2B00J+c2C00J+c2D00J+c2E00J+c2F00J;
assign A200J=(C200J>=0)?1:0;

assign P300J=A200J;

ninexnine_unit ninexnine_unit_5716(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2J000),
				.b1(W2J010),
				.b2(W2J020),
				.b3(W2J100),
				.b4(W2J110),
				.b5(W2J120),
				.b6(W2J200),
				.b7(W2J210),
				.b8(W2J220),
				.c(c2001J)
);

ninexnine_unit ninexnine_unit_5717(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2J001),
				.b1(W2J011),
				.b2(W2J021),
				.b3(W2J101),
				.b4(W2J111),
				.b5(W2J121),
				.b6(W2J201),
				.b7(W2J211),
				.b8(W2J221),
				.c(c2101J)
);

ninexnine_unit ninexnine_unit_5718(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2J002),
				.b1(W2J012),
				.b2(W2J022),
				.b3(W2J102),
				.b4(W2J112),
				.b5(W2J122),
				.b6(W2J202),
				.b7(W2J212),
				.b8(W2J222),
				.c(c2201J)
);

ninexnine_unit ninexnine_unit_5719(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2J003),
				.b1(W2J013),
				.b2(W2J023),
				.b3(W2J103),
				.b4(W2J113),
				.b5(W2J123),
				.b6(W2J203),
				.b7(W2J213),
				.b8(W2J223),
				.c(c2301J)
);

ninexnine_unit ninexnine_unit_5720(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2J004),
				.b1(W2J014),
				.b2(W2J024),
				.b3(W2J104),
				.b4(W2J114),
				.b5(W2J124),
				.b6(W2J204),
				.b7(W2J214),
				.b8(W2J224),
				.c(c2401J)
);

ninexnine_unit ninexnine_unit_5721(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2J005),
				.b1(W2J015),
				.b2(W2J025),
				.b3(W2J105),
				.b4(W2J115),
				.b5(W2J125),
				.b6(W2J205),
				.b7(W2J215),
				.b8(W2J225),
				.c(c2501J)
);

ninexnine_unit ninexnine_unit_5722(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2J006),
				.b1(W2J016),
				.b2(W2J026),
				.b3(W2J106),
				.b4(W2J116),
				.b5(W2J126),
				.b6(W2J206),
				.b7(W2J216),
				.b8(W2J226),
				.c(c2601J)
);

ninexnine_unit ninexnine_unit_5723(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2J007),
				.b1(W2J017),
				.b2(W2J027),
				.b3(W2J107),
				.b4(W2J117),
				.b5(W2J127),
				.b6(W2J207),
				.b7(W2J217),
				.b8(W2J227),
				.c(c2701J)
);

ninexnine_unit ninexnine_unit_5724(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2J008),
				.b1(W2J018),
				.b2(W2J028),
				.b3(W2J108),
				.b4(W2J118),
				.b5(W2J128),
				.b6(W2J208),
				.b7(W2J218),
				.b8(W2J228),
				.c(c2801J)
);

ninexnine_unit ninexnine_unit_5725(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2J009),
				.b1(W2J019),
				.b2(W2J029),
				.b3(W2J109),
				.b4(W2J119),
				.b5(W2J129),
				.b6(W2J209),
				.b7(W2J219),
				.b8(W2J229),
				.c(c2901J)
);

ninexnine_unit ninexnine_unit_5726(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2J00A),
				.b1(W2J01A),
				.b2(W2J02A),
				.b3(W2J10A),
				.b4(W2J11A),
				.b5(W2J12A),
				.b6(W2J20A),
				.b7(W2J21A),
				.b8(W2J22A),
				.c(c2A01J)
);

ninexnine_unit ninexnine_unit_5727(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2J00B),
				.b1(W2J01B),
				.b2(W2J02B),
				.b3(W2J10B),
				.b4(W2J11B),
				.b5(W2J12B),
				.b6(W2J20B),
				.b7(W2J21B),
				.b8(W2J22B),
				.c(c2B01J)
);

ninexnine_unit ninexnine_unit_5728(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2J00C),
				.b1(W2J01C),
				.b2(W2J02C),
				.b3(W2J10C),
				.b4(W2J11C),
				.b5(W2J12C),
				.b6(W2J20C),
				.b7(W2J21C),
				.b8(W2J22C),
				.c(c2C01J)
);

ninexnine_unit ninexnine_unit_5729(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2J00D),
				.b1(W2J01D),
				.b2(W2J02D),
				.b3(W2J10D),
				.b4(W2J11D),
				.b5(W2J12D),
				.b6(W2J20D),
				.b7(W2J21D),
				.b8(W2J22D),
				.c(c2D01J)
);

ninexnine_unit ninexnine_unit_5730(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2J00E),
				.b1(W2J01E),
				.b2(W2J02E),
				.b3(W2J10E),
				.b4(W2J11E),
				.b5(W2J12E),
				.b6(W2J20E),
				.b7(W2J21E),
				.b8(W2J22E),
				.c(c2E01J)
);

ninexnine_unit ninexnine_unit_5731(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2J00F),
				.b1(W2J01F),
				.b2(W2J02F),
				.b3(W2J10F),
				.b4(W2J11F),
				.b5(W2J12F),
				.b6(W2J20F),
				.b7(W2J21F),
				.b8(W2J22F),
				.c(c2F01J)
);

assign C201J=c2001J+c2101J+c2201J+c2301J+c2401J+c2501J+c2601J+c2701J+c2801J+c2901J+c2A01J+c2B01J+c2C01J+c2D01J+c2E01J+c2F01J;
assign A201J=(C201J>=0)?1:0;

assign P301J=A201J;

ninexnine_unit ninexnine_unit_5732(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2J000),
				.b1(W2J010),
				.b2(W2J020),
				.b3(W2J100),
				.b4(W2J110),
				.b5(W2J120),
				.b6(W2J200),
				.b7(W2J210),
				.b8(W2J220),
				.c(c2002J)
);

ninexnine_unit ninexnine_unit_5733(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2J001),
				.b1(W2J011),
				.b2(W2J021),
				.b3(W2J101),
				.b4(W2J111),
				.b5(W2J121),
				.b6(W2J201),
				.b7(W2J211),
				.b8(W2J221),
				.c(c2102J)
);

ninexnine_unit ninexnine_unit_5734(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2J002),
				.b1(W2J012),
				.b2(W2J022),
				.b3(W2J102),
				.b4(W2J112),
				.b5(W2J122),
				.b6(W2J202),
				.b7(W2J212),
				.b8(W2J222),
				.c(c2202J)
);

ninexnine_unit ninexnine_unit_5735(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2J003),
				.b1(W2J013),
				.b2(W2J023),
				.b3(W2J103),
				.b4(W2J113),
				.b5(W2J123),
				.b6(W2J203),
				.b7(W2J213),
				.b8(W2J223),
				.c(c2302J)
);

ninexnine_unit ninexnine_unit_5736(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2J004),
				.b1(W2J014),
				.b2(W2J024),
				.b3(W2J104),
				.b4(W2J114),
				.b5(W2J124),
				.b6(W2J204),
				.b7(W2J214),
				.b8(W2J224),
				.c(c2402J)
);

ninexnine_unit ninexnine_unit_5737(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2J005),
				.b1(W2J015),
				.b2(W2J025),
				.b3(W2J105),
				.b4(W2J115),
				.b5(W2J125),
				.b6(W2J205),
				.b7(W2J215),
				.b8(W2J225),
				.c(c2502J)
);

ninexnine_unit ninexnine_unit_5738(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2J006),
				.b1(W2J016),
				.b2(W2J026),
				.b3(W2J106),
				.b4(W2J116),
				.b5(W2J126),
				.b6(W2J206),
				.b7(W2J216),
				.b8(W2J226),
				.c(c2602J)
);

ninexnine_unit ninexnine_unit_5739(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2J007),
				.b1(W2J017),
				.b2(W2J027),
				.b3(W2J107),
				.b4(W2J117),
				.b5(W2J127),
				.b6(W2J207),
				.b7(W2J217),
				.b8(W2J227),
				.c(c2702J)
);

ninexnine_unit ninexnine_unit_5740(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2J008),
				.b1(W2J018),
				.b2(W2J028),
				.b3(W2J108),
				.b4(W2J118),
				.b5(W2J128),
				.b6(W2J208),
				.b7(W2J218),
				.b8(W2J228),
				.c(c2802J)
);

ninexnine_unit ninexnine_unit_5741(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2J009),
				.b1(W2J019),
				.b2(W2J029),
				.b3(W2J109),
				.b4(W2J119),
				.b5(W2J129),
				.b6(W2J209),
				.b7(W2J219),
				.b8(W2J229),
				.c(c2902J)
);

ninexnine_unit ninexnine_unit_5742(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2J00A),
				.b1(W2J01A),
				.b2(W2J02A),
				.b3(W2J10A),
				.b4(W2J11A),
				.b5(W2J12A),
				.b6(W2J20A),
				.b7(W2J21A),
				.b8(W2J22A),
				.c(c2A02J)
);

ninexnine_unit ninexnine_unit_5743(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2J00B),
				.b1(W2J01B),
				.b2(W2J02B),
				.b3(W2J10B),
				.b4(W2J11B),
				.b5(W2J12B),
				.b6(W2J20B),
				.b7(W2J21B),
				.b8(W2J22B),
				.c(c2B02J)
);

ninexnine_unit ninexnine_unit_5744(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2J00C),
				.b1(W2J01C),
				.b2(W2J02C),
				.b3(W2J10C),
				.b4(W2J11C),
				.b5(W2J12C),
				.b6(W2J20C),
				.b7(W2J21C),
				.b8(W2J22C),
				.c(c2C02J)
);

ninexnine_unit ninexnine_unit_5745(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2J00D),
				.b1(W2J01D),
				.b2(W2J02D),
				.b3(W2J10D),
				.b4(W2J11D),
				.b5(W2J12D),
				.b6(W2J20D),
				.b7(W2J21D),
				.b8(W2J22D),
				.c(c2D02J)
);

ninexnine_unit ninexnine_unit_5746(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2J00E),
				.b1(W2J01E),
				.b2(W2J02E),
				.b3(W2J10E),
				.b4(W2J11E),
				.b5(W2J12E),
				.b6(W2J20E),
				.b7(W2J21E),
				.b8(W2J22E),
				.c(c2E02J)
);

ninexnine_unit ninexnine_unit_5747(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2J00F),
				.b1(W2J01F),
				.b2(W2J02F),
				.b3(W2J10F),
				.b4(W2J11F),
				.b5(W2J12F),
				.b6(W2J20F),
				.b7(W2J21F),
				.b8(W2J22F),
				.c(c2F02J)
);

assign C202J=c2002J+c2102J+c2202J+c2302J+c2402J+c2502J+c2602J+c2702J+c2802J+c2902J+c2A02J+c2B02J+c2C02J+c2D02J+c2E02J+c2F02J;
assign A202J=(C202J>=0)?1:0;

assign P302J=A202J;

ninexnine_unit ninexnine_unit_5748(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2J000),
				.b1(W2J010),
				.b2(W2J020),
				.b3(W2J100),
				.b4(W2J110),
				.b5(W2J120),
				.b6(W2J200),
				.b7(W2J210),
				.b8(W2J220),
				.c(c2010J)
);

ninexnine_unit ninexnine_unit_5749(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2J001),
				.b1(W2J011),
				.b2(W2J021),
				.b3(W2J101),
				.b4(W2J111),
				.b5(W2J121),
				.b6(W2J201),
				.b7(W2J211),
				.b8(W2J221),
				.c(c2110J)
);

ninexnine_unit ninexnine_unit_5750(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2J002),
				.b1(W2J012),
				.b2(W2J022),
				.b3(W2J102),
				.b4(W2J112),
				.b5(W2J122),
				.b6(W2J202),
				.b7(W2J212),
				.b8(W2J222),
				.c(c2210J)
);

ninexnine_unit ninexnine_unit_5751(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2J003),
				.b1(W2J013),
				.b2(W2J023),
				.b3(W2J103),
				.b4(W2J113),
				.b5(W2J123),
				.b6(W2J203),
				.b7(W2J213),
				.b8(W2J223),
				.c(c2310J)
);

ninexnine_unit ninexnine_unit_5752(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2J004),
				.b1(W2J014),
				.b2(W2J024),
				.b3(W2J104),
				.b4(W2J114),
				.b5(W2J124),
				.b6(W2J204),
				.b7(W2J214),
				.b8(W2J224),
				.c(c2410J)
);

ninexnine_unit ninexnine_unit_5753(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2J005),
				.b1(W2J015),
				.b2(W2J025),
				.b3(W2J105),
				.b4(W2J115),
				.b5(W2J125),
				.b6(W2J205),
				.b7(W2J215),
				.b8(W2J225),
				.c(c2510J)
);

ninexnine_unit ninexnine_unit_5754(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2J006),
				.b1(W2J016),
				.b2(W2J026),
				.b3(W2J106),
				.b4(W2J116),
				.b5(W2J126),
				.b6(W2J206),
				.b7(W2J216),
				.b8(W2J226),
				.c(c2610J)
);

ninexnine_unit ninexnine_unit_5755(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2J007),
				.b1(W2J017),
				.b2(W2J027),
				.b3(W2J107),
				.b4(W2J117),
				.b5(W2J127),
				.b6(W2J207),
				.b7(W2J217),
				.b8(W2J227),
				.c(c2710J)
);

ninexnine_unit ninexnine_unit_5756(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2J008),
				.b1(W2J018),
				.b2(W2J028),
				.b3(W2J108),
				.b4(W2J118),
				.b5(W2J128),
				.b6(W2J208),
				.b7(W2J218),
				.b8(W2J228),
				.c(c2810J)
);

ninexnine_unit ninexnine_unit_5757(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2J009),
				.b1(W2J019),
				.b2(W2J029),
				.b3(W2J109),
				.b4(W2J119),
				.b5(W2J129),
				.b6(W2J209),
				.b7(W2J219),
				.b8(W2J229),
				.c(c2910J)
);

ninexnine_unit ninexnine_unit_5758(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2J00A),
				.b1(W2J01A),
				.b2(W2J02A),
				.b3(W2J10A),
				.b4(W2J11A),
				.b5(W2J12A),
				.b6(W2J20A),
				.b7(W2J21A),
				.b8(W2J22A),
				.c(c2A10J)
);

ninexnine_unit ninexnine_unit_5759(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2J00B),
				.b1(W2J01B),
				.b2(W2J02B),
				.b3(W2J10B),
				.b4(W2J11B),
				.b5(W2J12B),
				.b6(W2J20B),
				.b7(W2J21B),
				.b8(W2J22B),
				.c(c2B10J)
);

ninexnine_unit ninexnine_unit_5760(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2J00C),
				.b1(W2J01C),
				.b2(W2J02C),
				.b3(W2J10C),
				.b4(W2J11C),
				.b5(W2J12C),
				.b6(W2J20C),
				.b7(W2J21C),
				.b8(W2J22C),
				.c(c2C10J)
);

ninexnine_unit ninexnine_unit_5761(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2J00D),
				.b1(W2J01D),
				.b2(W2J02D),
				.b3(W2J10D),
				.b4(W2J11D),
				.b5(W2J12D),
				.b6(W2J20D),
				.b7(W2J21D),
				.b8(W2J22D),
				.c(c2D10J)
);

ninexnine_unit ninexnine_unit_5762(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2J00E),
				.b1(W2J01E),
				.b2(W2J02E),
				.b3(W2J10E),
				.b4(W2J11E),
				.b5(W2J12E),
				.b6(W2J20E),
				.b7(W2J21E),
				.b8(W2J22E),
				.c(c2E10J)
);

ninexnine_unit ninexnine_unit_5763(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2J00F),
				.b1(W2J01F),
				.b2(W2J02F),
				.b3(W2J10F),
				.b4(W2J11F),
				.b5(W2J12F),
				.b6(W2J20F),
				.b7(W2J21F),
				.b8(W2J22F),
				.c(c2F10J)
);

assign C210J=c2010J+c2110J+c2210J+c2310J+c2410J+c2510J+c2610J+c2710J+c2810J+c2910J+c2A10J+c2B10J+c2C10J+c2D10J+c2E10J+c2F10J;
assign A210J=(C210J>=0)?1:0;

assign P310J=A210J;

ninexnine_unit ninexnine_unit_5764(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2J000),
				.b1(W2J010),
				.b2(W2J020),
				.b3(W2J100),
				.b4(W2J110),
				.b5(W2J120),
				.b6(W2J200),
				.b7(W2J210),
				.b8(W2J220),
				.c(c2011J)
);

ninexnine_unit ninexnine_unit_5765(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2J001),
				.b1(W2J011),
				.b2(W2J021),
				.b3(W2J101),
				.b4(W2J111),
				.b5(W2J121),
				.b6(W2J201),
				.b7(W2J211),
				.b8(W2J221),
				.c(c2111J)
);

ninexnine_unit ninexnine_unit_5766(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2J002),
				.b1(W2J012),
				.b2(W2J022),
				.b3(W2J102),
				.b4(W2J112),
				.b5(W2J122),
				.b6(W2J202),
				.b7(W2J212),
				.b8(W2J222),
				.c(c2211J)
);

ninexnine_unit ninexnine_unit_5767(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2J003),
				.b1(W2J013),
				.b2(W2J023),
				.b3(W2J103),
				.b4(W2J113),
				.b5(W2J123),
				.b6(W2J203),
				.b7(W2J213),
				.b8(W2J223),
				.c(c2311J)
);

ninexnine_unit ninexnine_unit_5768(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2J004),
				.b1(W2J014),
				.b2(W2J024),
				.b3(W2J104),
				.b4(W2J114),
				.b5(W2J124),
				.b6(W2J204),
				.b7(W2J214),
				.b8(W2J224),
				.c(c2411J)
);

ninexnine_unit ninexnine_unit_5769(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2J005),
				.b1(W2J015),
				.b2(W2J025),
				.b3(W2J105),
				.b4(W2J115),
				.b5(W2J125),
				.b6(W2J205),
				.b7(W2J215),
				.b8(W2J225),
				.c(c2511J)
);

ninexnine_unit ninexnine_unit_5770(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2J006),
				.b1(W2J016),
				.b2(W2J026),
				.b3(W2J106),
				.b4(W2J116),
				.b5(W2J126),
				.b6(W2J206),
				.b7(W2J216),
				.b8(W2J226),
				.c(c2611J)
);

ninexnine_unit ninexnine_unit_5771(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2J007),
				.b1(W2J017),
				.b2(W2J027),
				.b3(W2J107),
				.b4(W2J117),
				.b5(W2J127),
				.b6(W2J207),
				.b7(W2J217),
				.b8(W2J227),
				.c(c2711J)
);

ninexnine_unit ninexnine_unit_5772(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2J008),
				.b1(W2J018),
				.b2(W2J028),
				.b3(W2J108),
				.b4(W2J118),
				.b5(W2J128),
				.b6(W2J208),
				.b7(W2J218),
				.b8(W2J228),
				.c(c2811J)
);

ninexnine_unit ninexnine_unit_5773(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2J009),
				.b1(W2J019),
				.b2(W2J029),
				.b3(W2J109),
				.b4(W2J119),
				.b5(W2J129),
				.b6(W2J209),
				.b7(W2J219),
				.b8(W2J229),
				.c(c2911J)
);

ninexnine_unit ninexnine_unit_5774(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2J00A),
				.b1(W2J01A),
				.b2(W2J02A),
				.b3(W2J10A),
				.b4(W2J11A),
				.b5(W2J12A),
				.b6(W2J20A),
				.b7(W2J21A),
				.b8(W2J22A),
				.c(c2A11J)
);

ninexnine_unit ninexnine_unit_5775(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2J00B),
				.b1(W2J01B),
				.b2(W2J02B),
				.b3(W2J10B),
				.b4(W2J11B),
				.b5(W2J12B),
				.b6(W2J20B),
				.b7(W2J21B),
				.b8(W2J22B),
				.c(c2B11J)
);

ninexnine_unit ninexnine_unit_5776(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2J00C),
				.b1(W2J01C),
				.b2(W2J02C),
				.b3(W2J10C),
				.b4(W2J11C),
				.b5(W2J12C),
				.b6(W2J20C),
				.b7(W2J21C),
				.b8(W2J22C),
				.c(c2C11J)
);

ninexnine_unit ninexnine_unit_5777(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2J00D),
				.b1(W2J01D),
				.b2(W2J02D),
				.b3(W2J10D),
				.b4(W2J11D),
				.b5(W2J12D),
				.b6(W2J20D),
				.b7(W2J21D),
				.b8(W2J22D),
				.c(c2D11J)
);

ninexnine_unit ninexnine_unit_5778(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2J00E),
				.b1(W2J01E),
				.b2(W2J02E),
				.b3(W2J10E),
				.b4(W2J11E),
				.b5(W2J12E),
				.b6(W2J20E),
				.b7(W2J21E),
				.b8(W2J22E),
				.c(c2E11J)
);

ninexnine_unit ninexnine_unit_5779(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2J00F),
				.b1(W2J01F),
				.b2(W2J02F),
				.b3(W2J10F),
				.b4(W2J11F),
				.b5(W2J12F),
				.b6(W2J20F),
				.b7(W2J21F),
				.b8(W2J22F),
				.c(c2F11J)
);

assign C211J=c2011J+c2111J+c2211J+c2311J+c2411J+c2511J+c2611J+c2711J+c2811J+c2911J+c2A11J+c2B11J+c2C11J+c2D11J+c2E11J+c2F11J;
assign A211J=(C211J>=0)?1:0;

assign P311J=A211J;

ninexnine_unit ninexnine_unit_5780(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2J000),
				.b1(W2J010),
				.b2(W2J020),
				.b3(W2J100),
				.b4(W2J110),
				.b5(W2J120),
				.b6(W2J200),
				.b7(W2J210),
				.b8(W2J220),
				.c(c2012J)
);

ninexnine_unit ninexnine_unit_5781(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2J001),
				.b1(W2J011),
				.b2(W2J021),
				.b3(W2J101),
				.b4(W2J111),
				.b5(W2J121),
				.b6(W2J201),
				.b7(W2J211),
				.b8(W2J221),
				.c(c2112J)
);

ninexnine_unit ninexnine_unit_5782(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2J002),
				.b1(W2J012),
				.b2(W2J022),
				.b3(W2J102),
				.b4(W2J112),
				.b5(W2J122),
				.b6(W2J202),
				.b7(W2J212),
				.b8(W2J222),
				.c(c2212J)
);

ninexnine_unit ninexnine_unit_5783(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2J003),
				.b1(W2J013),
				.b2(W2J023),
				.b3(W2J103),
				.b4(W2J113),
				.b5(W2J123),
				.b6(W2J203),
				.b7(W2J213),
				.b8(W2J223),
				.c(c2312J)
);

ninexnine_unit ninexnine_unit_5784(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2J004),
				.b1(W2J014),
				.b2(W2J024),
				.b3(W2J104),
				.b4(W2J114),
				.b5(W2J124),
				.b6(W2J204),
				.b7(W2J214),
				.b8(W2J224),
				.c(c2412J)
);

ninexnine_unit ninexnine_unit_5785(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2J005),
				.b1(W2J015),
				.b2(W2J025),
				.b3(W2J105),
				.b4(W2J115),
				.b5(W2J125),
				.b6(W2J205),
				.b7(W2J215),
				.b8(W2J225),
				.c(c2512J)
);

ninexnine_unit ninexnine_unit_5786(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2J006),
				.b1(W2J016),
				.b2(W2J026),
				.b3(W2J106),
				.b4(W2J116),
				.b5(W2J126),
				.b6(W2J206),
				.b7(W2J216),
				.b8(W2J226),
				.c(c2612J)
);

ninexnine_unit ninexnine_unit_5787(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2J007),
				.b1(W2J017),
				.b2(W2J027),
				.b3(W2J107),
				.b4(W2J117),
				.b5(W2J127),
				.b6(W2J207),
				.b7(W2J217),
				.b8(W2J227),
				.c(c2712J)
);

ninexnine_unit ninexnine_unit_5788(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2J008),
				.b1(W2J018),
				.b2(W2J028),
				.b3(W2J108),
				.b4(W2J118),
				.b5(W2J128),
				.b6(W2J208),
				.b7(W2J218),
				.b8(W2J228),
				.c(c2812J)
);

ninexnine_unit ninexnine_unit_5789(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2J009),
				.b1(W2J019),
				.b2(W2J029),
				.b3(W2J109),
				.b4(W2J119),
				.b5(W2J129),
				.b6(W2J209),
				.b7(W2J219),
				.b8(W2J229),
				.c(c2912J)
);

ninexnine_unit ninexnine_unit_5790(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2J00A),
				.b1(W2J01A),
				.b2(W2J02A),
				.b3(W2J10A),
				.b4(W2J11A),
				.b5(W2J12A),
				.b6(W2J20A),
				.b7(W2J21A),
				.b8(W2J22A),
				.c(c2A12J)
);

ninexnine_unit ninexnine_unit_5791(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2J00B),
				.b1(W2J01B),
				.b2(W2J02B),
				.b3(W2J10B),
				.b4(W2J11B),
				.b5(W2J12B),
				.b6(W2J20B),
				.b7(W2J21B),
				.b8(W2J22B),
				.c(c2B12J)
);

ninexnine_unit ninexnine_unit_5792(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2J00C),
				.b1(W2J01C),
				.b2(W2J02C),
				.b3(W2J10C),
				.b4(W2J11C),
				.b5(W2J12C),
				.b6(W2J20C),
				.b7(W2J21C),
				.b8(W2J22C),
				.c(c2C12J)
);

ninexnine_unit ninexnine_unit_5793(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2J00D),
				.b1(W2J01D),
				.b2(W2J02D),
				.b3(W2J10D),
				.b4(W2J11D),
				.b5(W2J12D),
				.b6(W2J20D),
				.b7(W2J21D),
				.b8(W2J22D),
				.c(c2D12J)
);

ninexnine_unit ninexnine_unit_5794(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2J00E),
				.b1(W2J01E),
				.b2(W2J02E),
				.b3(W2J10E),
				.b4(W2J11E),
				.b5(W2J12E),
				.b6(W2J20E),
				.b7(W2J21E),
				.b8(W2J22E),
				.c(c2E12J)
);

ninexnine_unit ninexnine_unit_5795(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2J00F),
				.b1(W2J01F),
				.b2(W2J02F),
				.b3(W2J10F),
				.b4(W2J11F),
				.b5(W2J12F),
				.b6(W2J20F),
				.b7(W2J21F),
				.b8(W2J22F),
				.c(c2F12J)
);

assign C212J=c2012J+c2112J+c2212J+c2312J+c2412J+c2512J+c2612J+c2712J+c2812J+c2912J+c2A12J+c2B12J+c2C12J+c2D12J+c2E12J+c2F12J;
assign A212J=(C212J>=0)?1:0;

assign P312J=A212J;

ninexnine_unit ninexnine_unit_5796(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2J000),
				.b1(W2J010),
				.b2(W2J020),
				.b3(W2J100),
				.b4(W2J110),
				.b5(W2J120),
				.b6(W2J200),
				.b7(W2J210),
				.b8(W2J220),
				.c(c2020J)
);

ninexnine_unit ninexnine_unit_5797(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2J001),
				.b1(W2J011),
				.b2(W2J021),
				.b3(W2J101),
				.b4(W2J111),
				.b5(W2J121),
				.b6(W2J201),
				.b7(W2J211),
				.b8(W2J221),
				.c(c2120J)
);

ninexnine_unit ninexnine_unit_5798(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2J002),
				.b1(W2J012),
				.b2(W2J022),
				.b3(W2J102),
				.b4(W2J112),
				.b5(W2J122),
				.b6(W2J202),
				.b7(W2J212),
				.b8(W2J222),
				.c(c2220J)
);

ninexnine_unit ninexnine_unit_5799(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2J003),
				.b1(W2J013),
				.b2(W2J023),
				.b3(W2J103),
				.b4(W2J113),
				.b5(W2J123),
				.b6(W2J203),
				.b7(W2J213),
				.b8(W2J223),
				.c(c2320J)
);

ninexnine_unit ninexnine_unit_5800(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2J004),
				.b1(W2J014),
				.b2(W2J024),
				.b3(W2J104),
				.b4(W2J114),
				.b5(W2J124),
				.b6(W2J204),
				.b7(W2J214),
				.b8(W2J224),
				.c(c2420J)
);

ninexnine_unit ninexnine_unit_5801(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2J005),
				.b1(W2J015),
				.b2(W2J025),
				.b3(W2J105),
				.b4(W2J115),
				.b5(W2J125),
				.b6(W2J205),
				.b7(W2J215),
				.b8(W2J225),
				.c(c2520J)
);

ninexnine_unit ninexnine_unit_5802(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2J006),
				.b1(W2J016),
				.b2(W2J026),
				.b3(W2J106),
				.b4(W2J116),
				.b5(W2J126),
				.b6(W2J206),
				.b7(W2J216),
				.b8(W2J226),
				.c(c2620J)
);

ninexnine_unit ninexnine_unit_5803(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2J007),
				.b1(W2J017),
				.b2(W2J027),
				.b3(W2J107),
				.b4(W2J117),
				.b5(W2J127),
				.b6(W2J207),
				.b7(W2J217),
				.b8(W2J227),
				.c(c2720J)
);

ninexnine_unit ninexnine_unit_5804(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2J008),
				.b1(W2J018),
				.b2(W2J028),
				.b3(W2J108),
				.b4(W2J118),
				.b5(W2J128),
				.b6(W2J208),
				.b7(W2J218),
				.b8(W2J228),
				.c(c2820J)
);

ninexnine_unit ninexnine_unit_5805(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2J009),
				.b1(W2J019),
				.b2(W2J029),
				.b3(W2J109),
				.b4(W2J119),
				.b5(W2J129),
				.b6(W2J209),
				.b7(W2J219),
				.b8(W2J229),
				.c(c2920J)
);

ninexnine_unit ninexnine_unit_5806(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2J00A),
				.b1(W2J01A),
				.b2(W2J02A),
				.b3(W2J10A),
				.b4(W2J11A),
				.b5(W2J12A),
				.b6(W2J20A),
				.b7(W2J21A),
				.b8(W2J22A),
				.c(c2A20J)
);

ninexnine_unit ninexnine_unit_5807(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2J00B),
				.b1(W2J01B),
				.b2(W2J02B),
				.b3(W2J10B),
				.b4(W2J11B),
				.b5(W2J12B),
				.b6(W2J20B),
				.b7(W2J21B),
				.b8(W2J22B),
				.c(c2B20J)
);

ninexnine_unit ninexnine_unit_5808(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2J00C),
				.b1(W2J01C),
				.b2(W2J02C),
				.b3(W2J10C),
				.b4(W2J11C),
				.b5(W2J12C),
				.b6(W2J20C),
				.b7(W2J21C),
				.b8(W2J22C),
				.c(c2C20J)
);

ninexnine_unit ninexnine_unit_5809(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2J00D),
				.b1(W2J01D),
				.b2(W2J02D),
				.b3(W2J10D),
				.b4(W2J11D),
				.b5(W2J12D),
				.b6(W2J20D),
				.b7(W2J21D),
				.b8(W2J22D),
				.c(c2D20J)
);

ninexnine_unit ninexnine_unit_5810(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2J00E),
				.b1(W2J01E),
				.b2(W2J02E),
				.b3(W2J10E),
				.b4(W2J11E),
				.b5(W2J12E),
				.b6(W2J20E),
				.b7(W2J21E),
				.b8(W2J22E),
				.c(c2E20J)
);

ninexnine_unit ninexnine_unit_5811(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2J00F),
				.b1(W2J01F),
				.b2(W2J02F),
				.b3(W2J10F),
				.b4(W2J11F),
				.b5(W2J12F),
				.b6(W2J20F),
				.b7(W2J21F),
				.b8(W2J22F),
				.c(c2F20J)
);

assign C220J=c2020J+c2120J+c2220J+c2320J+c2420J+c2520J+c2620J+c2720J+c2820J+c2920J+c2A20J+c2B20J+c2C20J+c2D20J+c2E20J+c2F20J;
assign A220J=(C220J>=0)?1:0;

assign P320J=A220J;

ninexnine_unit ninexnine_unit_5812(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2J000),
				.b1(W2J010),
				.b2(W2J020),
				.b3(W2J100),
				.b4(W2J110),
				.b5(W2J120),
				.b6(W2J200),
				.b7(W2J210),
				.b8(W2J220),
				.c(c2021J)
);

ninexnine_unit ninexnine_unit_5813(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2J001),
				.b1(W2J011),
				.b2(W2J021),
				.b3(W2J101),
				.b4(W2J111),
				.b5(W2J121),
				.b6(W2J201),
				.b7(W2J211),
				.b8(W2J221),
				.c(c2121J)
);

ninexnine_unit ninexnine_unit_5814(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2J002),
				.b1(W2J012),
				.b2(W2J022),
				.b3(W2J102),
				.b4(W2J112),
				.b5(W2J122),
				.b6(W2J202),
				.b7(W2J212),
				.b8(W2J222),
				.c(c2221J)
);

ninexnine_unit ninexnine_unit_5815(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2J003),
				.b1(W2J013),
				.b2(W2J023),
				.b3(W2J103),
				.b4(W2J113),
				.b5(W2J123),
				.b6(W2J203),
				.b7(W2J213),
				.b8(W2J223),
				.c(c2321J)
);

ninexnine_unit ninexnine_unit_5816(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2J004),
				.b1(W2J014),
				.b2(W2J024),
				.b3(W2J104),
				.b4(W2J114),
				.b5(W2J124),
				.b6(W2J204),
				.b7(W2J214),
				.b8(W2J224),
				.c(c2421J)
);

ninexnine_unit ninexnine_unit_5817(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2J005),
				.b1(W2J015),
				.b2(W2J025),
				.b3(W2J105),
				.b4(W2J115),
				.b5(W2J125),
				.b6(W2J205),
				.b7(W2J215),
				.b8(W2J225),
				.c(c2521J)
);

ninexnine_unit ninexnine_unit_5818(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2J006),
				.b1(W2J016),
				.b2(W2J026),
				.b3(W2J106),
				.b4(W2J116),
				.b5(W2J126),
				.b6(W2J206),
				.b7(W2J216),
				.b8(W2J226),
				.c(c2621J)
);

ninexnine_unit ninexnine_unit_5819(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2J007),
				.b1(W2J017),
				.b2(W2J027),
				.b3(W2J107),
				.b4(W2J117),
				.b5(W2J127),
				.b6(W2J207),
				.b7(W2J217),
				.b8(W2J227),
				.c(c2721J)
);

ninexnine_unit ninexnine_unit_5820(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2J008),
				.b1(W2J018),
				.b2(W2J028),
				.b3(W2J108),
				.b4(W2J118),
				.b5(W2J128),
				.b6(W2J208),
				.b7(W2J218),
				.b8(W2J228),
				.c(c2821J)
);

ninexnine_unit ninexnine_unit_5821(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2J009),
				.b1(W2J019),
				.b2(W2J029),
				.b3(W2J109),
				.b4(W2J119),
				.b5(W2J129),
				.b6(W2J209),
				.b7(W2J219),
				.b8(W2J229),
				.c(c2921J)
);

ninexnine_unit ninexnine_unit_5822(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2J00A),
				.b1(W2J01A),
				.b2(W2J02A),
				.b3(W2J10A),
				.b4(W2J11A),
				.b5(W2J12A),
				.b6(W2J20A),
				.b7(W2J21A),
				.b8(W2J22A),
				.c(c2A21J)
);

ninexnine_unit ninexnine_unit_5823(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2J00B),
				.b1(W2J01B),
				.b2(W2J02B),
				.b3(W2J10B),
				.b4(W2J11B),
				.b5(W2J12B),
				.b6(W2J20B),
				.b7(W2J21B),
				.b8(W2J22B),
				.c(c2B21J)
);

ninexnine_unit ninexnine_unit_5824(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2J00C),
				.b1(W2J01C),
				.b2(W2J02C),
				.b3(W2J10C),
				.b4(W2J11C),
				.b5(W2J12C),
				.b6(W2J20C),
				.b7(W2J21C),
				.b8(W2J22C),
				.c(c2C21J)
);

ninexnine_unit ninexnine_unit_5825(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2J00D),
				.b1(W2J01D),
				.b2(W2J02D),
				.b3(W2J10D),
				.b4(W2J11D),
				.b5(W2J12D),
				.b6(W2J20D),
				.b7(W2J21D),
				.b8(W2J22D),
				.c(c2D21J)
);

ninexnine_unit ninexnine_unit_5826(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2J00E),
				.b1(W2J01E),
				.b2(W2J02E),
				.b3(W2J10E),
				.b4(W2J11E),
				.b5(W2J12E),
				.b6(W2J20E),
				.b7(W2J21E),
				.b8(W2J22E),
				.c(c2E21J)
);

ninexnine_unit ninexnine_unit_5827(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2J00F),
				.b1(W2J01F),
				.b2(W2J02F),
				.b3(W2J10F),
				.b4(W2J11F),
				.b5(W2J12F),
				.b6(W2J20F),
				.b7(W2J21F),
				.b8(W2J22F),
				.c(c2F21J)
);

assign C221J=c2021J+c2121J+c2221J+c2321J+c2421J+c2521J+c2621J+c2721J+c2821J+c2921J+c2A21J+c2B21J+c2C21J+c2D21J+c2E21J+c2F21J;
assign A221J=(C221J>=0)?1:0;

assign P321J=A221J;

ninexnine_unit ninexnine_unit_5828(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2J000),
				.b1(W2J010),
				.b2(W2J020),
				.b3(W2J100),
				.b4(W2J110),
				.b5(W2J120),
				.b6(W2J200),
				.b7(W2J210),
				.b8(W2J220),
				.c(c2022J)
);

ninexnine_unit ninexnine_unit_5829(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2J001),
				.b1(W2J011),
				.b2(W2J021),
				.b3(W2J101),
				.b4(W2J111),
				.b5(W2J121),
				.b6(W2J201),
				.b7(W2J211),
				.b8(W2J221),
				.c(c2122J)
);

ninexnine_unit ninexnine_unit_5830(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2J002),
				.b1(W2J012),
				.b2(W2J022),
				.b3(W2J102),
				.b4(W2J112),
				.b5(W2J122),
				.b6(W2J202),
				.b7(W2J212),
				.b8(W2J222),
				.c(c2222J)
);

ninexnine_unit ninexnine_unit_5831(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2J003),
				.b1(W2J013),
				.b2(W2J023),
				.b3(W2J103),
				.b4(W2J113),
				.b5(W2J123),
				.b6(W2J203),
				.b7(W2J213),
				.b8(W2J223),
				.c(c2322J)
);

ninexnine_unit ninexnine_unit_5832(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2J004),
				.b1(W2J014),
				.b2(W2J024),
				.b3(W2J104),
				.b4(W2J114),
				.b5(W2J124),
				.b6(W2J204),
				.b7(W2J214),
				.b8(W2J224),
				.c(c2422J)
);

ninexnine_unit ninexnine_unit_5833(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2J005),
				.b1(W2J015),
				.b2(W2J025),
				.b3(W2J105),
				.b4(W2J115),
				.b5(W2J125),
				.b6(W2J205),
				.b7(W2J215),
				.b8(W2J225),
				.c(c2522J)
);

ninexnine_unit ninexnine_unit_5834(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2J006),
				.b1(W2J016),
				.b2(W2J026),
				.b3(W2J106),
				.b4(W2J116),
				.b5(W2J126),
				.b6(W2J206),
				.b7(W2J216),
				.b8(W2J226),
				.c(c2622J)
);

ninexnine_unit ninexnine_unit_5835(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2J007),
				.b1(W2J017),
				.b2(W2J027),
				.b3(W2J107),
				.b4(W2J117),
				.b5(W2J127),
				.b6(W2J207),
				.b7(W2J217),
				.b8(W2J227),
				.c(c2722J)
);

ninexnine_unit ninexnine_unit_5836(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2J008),
				.b1(W2J018),
				.b2(W2J028),
				.b3(W2J108),
				.b4(W2J118),
				.b5(W2J128),
				.b6(W2J208),
				.b7(W2J218),
				.b8(W2J228),
				.c(c2822J)
);

ninexnine_unit ninexnine_unit_5837(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2J009),
				.b1(W2J019),
				.b2(W2J029),
				.b3(W2J109),
				.b4(W2J119),
				.b5(W2J129),
				.b6(W2J209),
				.b7(W2J219),
				.b8(W2J229),
				.c(c2922J)
);

ninexnine_unit ninexnine_unit_5838(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2J00A),
				.b1(W2J01A),
				.b2(W2J02A),
				.b3(W2J10A),
				.b4(W2J11A),
				.b5(W2J12A),
				.b6(W2J20A),
				.b7(W2J21A),
				.b8(W2J22A),
				.c(c2A22J)
);

ninexnine_unit ninexnine_unit_5839(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2J00B),
				.b1(W2J01B),
				.b2(W2J02B),
				.b3(W2J10B),
				.b4(W2J11B),
				.b5(W2J12B),
				.b6(W2J20B),
				.b7(W2J21B),
				.b8(W2J22B),
				.c(c2B22J)
);

ninexnine_unit ninexnine_unit_5840(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2J00C),
				.b1(W2J01C),
				.b2(W2J02C),
				.b3(W2J10C),
				.b4(W2J11C),
				.b5(W2J12C),
				.b6(W2J20C),
				.b7(W2J21C),
				.b8(W2J22C),
				.c(c2C22J)
);

ninexnine_unit ninexnine_unit_5841(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2J00D),
				.b1(W2J01D),
				.b2(W2J02D),
				.b3(W2J10D),
				.b4(W2J11D),
				.b5(W2J12D),
				.b6(W2J20D),
				.b7(W2J21D),
				.b8(W2J22D),
				.c(c2D22J)
);

ninexnine_unit ninexnine_unit_5842(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2J00E),
				.b1(W2J01E),
				.b2(W2J02E),
				.b3(W2J10E),
				.b4(W2J11E),
				.b5(W2J12E),
				.b6(W2J20E),
				.b7(W2J21E),
				.b8(W2J22E),
				.c(c2E22J)
);

ninexnine_unit ninexnine_unit_5843(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2J00F),
				.b1(W2J01F),
				.b2(W2J02F),
				.b3(W2J10F),
				.b4(W2J11F),
				.b5(W2J12F),
				.b6(W2J20F),
				.b7(W2J21F),
				.b8(W2J22F),
				.c(c2F22J)
);

assign C222J=c2022J+c2122J+c2222J+c2322J+c2422J+c2522J+c2622J+c2722J+c2822J+c2922J+c2A22J+c2B22J+c2C22J+c2D22J+c2E22J+c2F22J;
assign A222J=(C222J>=0)?1:0;

assign P322J=A222J;

ninexnine_unit ninexnine_unit_5844(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2K000),
				.b1(W2K010),
				.b2(W2K020),
				.b3(W2K100),
				.b4(W2K110),
				.b5(W2K120),
				.b6(W2K200),
				.b7(W2K210),
				.b8(W2K220),
				.c(c2000K)
);

ninexnine_unit ninexnine_unit_5845(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2K001),
				.b1(W2K011),
				.b2(W2K021),
				.b3(W2K101),
				.b4(W2K111),
				.b5(W2K121),
				.b6(W2K201),
				.b7(W2K211),
				.b8(W2K221),
				.c(c2100K)
);

ninexnine_unit ninexnine_unit_5846(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2K002),
				.b1(W2K012),
				.b2(W2K022),
				.b3(W2K102),
				.b4(W2K112),
				.b5(W2K122),
				.b6(W2K202),
				.b7(W2K212),
				.b8(W2K222),
				.c(c2200K)
);

ninexnine_unit ninexnine_unit_5847(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2K003),
				.b1(W2K013),
				.b2(W2K023),
				.b3(W2K103),
				.b4(W2K113),
				.b5(W2K123),
				.b6(W2K203),
				.b7(W2K213),
				.b8(W2K223),
				.c(c2300K)
);

ninexnine_unit ninexnine_unit_5848(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2K004),
				.b1(W2K014),
				.b2(W2K024),
				.b3(W2K104),
				.b4(W2K114),
				.b5(W2K124),
				.b6(W2K204),
				.b7(W2K214),
				.b8(W2K224),
				.c(c2400K)
);

ninexnine_unit ninexnine_unit_5849(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2K005),
				.b1(W2K015),
				.b2(W2K025),
				.b3(W2K105),
				.b4(W2K115),
				.b5(W2K125),
				.b6(W2K205),
				.b7(W2K215),
				.b8(W2K225),
				.c(c2500K)
);

ninexnine_unit ninexnine_unit_5850(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2K006),
				.b1(W2K016),
				.b2(W2K026),
				.b3(W2K106),
				.b4(W2K116),
				.b5(W2K126),
				.b6(W2K206),
				.b7(W2K216),
				.b8(W2K226),
				.c(c2600K)
);

ninexnine_unit ninexnine_unit_5851(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2K007),
				.b1(W2K017),
				.b2(W2K027),
				.b3(W2K107),
				.b4(W2K117),
				.b5(W2K127),
				.b6(W2K207),
				.b7(W2K217),
				.b8(W2K227),
				.c(c2700K)
);

ninexnine_unit ninexnine_unit_5852(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2K008),
				.b1(W2K018),
				.b2(W2K028),
				.b3(W2K108),
				.b4(W2K118),
				.b5(W2K128),
				.b6(W2K208),
				.b7(W2K218),
				.b8(W2K228),
				.c(c2800K)
);

ninexnine_unit ninexnine_unit_5853(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2K009),
				.b1(W2K019),
				.b2(W2K029),
				.b3(W2K109),
				.b4(W2K119),
				.b5(W2K129),
				.b6(W2K209),
				.b7(W2K219),
				.b8(W2K229),
				.c(c2900K)
);

ninexnine_unit ninexnine_unit_5854(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2K00A),
				.b1(W2K01A),
				.b2(W2K02A),
				.b3(W2K10A),
				.b4(W2K11A),
				.b5(W2K12A),
				.b6(W2K20A),
				.b7(W2K21A),
				.b8(W2K22A),
				.c(c2A00K)
);

ninexnine_unit ninexnine_unit_5855(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2K00B),
				.b1(W2K01B),
				.b2(W2K02B),
				.b3(W2K10B),
				.b4(W2K11B),
				.b5(W2K12B),
				.b6(W2K20B),
				.b7(W2K21B),
				.b8(W2K22B),
				.c(c2B00K)
);

ninexnine_unit ninexnine_unit_5856(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2K00C),
				.b1(W2K01C),
				.b2(W2K02C),
				.b3(W2K10C),
				.b4(W2K11C),
				.b5(W2K12C),
				.b6(W2K20C),
				.b7(W2K21C),
				.b8(W2K22C),
				.c(c2C00K)
);

ninexnine_unit ninexnine_unit_5857(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2K00D),
				.b1(W2K01D),
				.b2(W2K02D),
				.b3(W2K10D),
				.b4(W2K11D),
				.b5(W2K12D),
				.b6(W2K20D),
				.b7(W2K21D),
				.b8(W2K22D),
				.c(c2D00K)
);

ninexnine_unit ninexnine_unit_5858(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2K00E),
				.b1(W2K01E),
				.b2(W2K02E),
				.b3(W2K10E),
				.b4(W2K11E),
				.b5(W2K12E),
				.b6(W2K20E),
				.b7(W2K21E),
				.b8(W2K22E),
				.c(c2E00K)
);

ninexnine_unit ninexnine_unit_5859(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2K00F),
				.b1(W2K01F),
				.b2(W2K02F),
				.b3(W2K10F),
				.b4(W2K11F),
				.b5(W2K12F),
				.b6(W2K20F),
				.b7(W2K21F),
				.b8(W2K22F),
				.c(c2F00K)
);

assign C200K=c2000K+c2100K+c2200K+c2300K+c2400K+c2500K+c2600K+c2700K+c2800K+c2900K+c2A00K+c2B00K+c2C00K+c2D00K+c2E00K+c2F00K;
assign A200K=(C200K>=0)?1:0;

assign P300K=A200K;

ninexnine_unit ninexnine_unit_5860(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2K000),
				.b1(W2K010),
				.b2(W2K020),
				.b3(W2K100),
				.b4(W2K110),
				.b5(W2K120),
				.b6(W2K200),
				.b7(W2K210),
				.b8(W2K220),
				.c(c2001K)
);

ninexnine_unit ninexnine_unit_5861(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2K001),
				.b1(W2K011),
				.b2(W2K021),
				.b3(W2K101),
				.b4(W2K111),
				.b5(W2K121),
				.b6(W2K201),
				.b7(W2K211),
				.b8(W2K221),
				.c(c2101K)
);

ninexnine_unit ninexnine_unit_5862(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2K002),
				.b1(W2K012),
				.b2(W2K022),
				.b3(W2K102),
				.b4(W2K112),
				.b5(W2K122),
				.b6(W2K202),
				.b7(W2K212),
				.b8(W2K222),
				.c(c2201K)
);

ninexnine_unit ninexnine_unit_5863(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2K003),
				.b1(W2K013),
				.b2(W2K023),
				.b3(W2K103),
				.b4(W2K113),
				.b5(W2K123),
				.b6(W2K203),
				.b7(W2K213),
				.b8(W2K223),
				.c(c2301K)
);

ninexnine_unit ninexnine_unit_5864(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2K004),
				.b1(W2K014),
				.b2(W2K024),
				.b3(W2K104),
				.b4(W2K114),
				.b5(W2K124),
				.b6(W2K204),
				.b7(W2K214),
				.b8(W2K224),
				.c(c2401K)
);

ninexnine_unit ninexnine_unit_5865(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2K005),
				.b1(W2K015),
				.b2(W2K025),
				.b3(W2K105),
				.b4(W2K115),
				.b5(W2K125),
				.b6(W2K205),
				.b7(W2K215),
				.b8(W2K225),
				.c(c2501K)
);

ninexnine_unit ninexnine_unit_5866(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2K006),
				.b1(W2K016),
				.b2(W2K026),
				.b3(W2K106),
				.b4(W2K116),
				.b5(W2K126),
				.b6(W2K206),
				.b7(W2K216),
				.b8(W2K226),
				.c(c2601K)
);

ninexnine_unit ninexnine_unit_5867(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2K007),
				.b1(W2K017),
				.b2(W2K027),
				.b3(W2K107),
				.b4(W2K117),
				.b5(W2K127),
				.b6(W2K207),
				.b7(W2K217),
				.b8(W2K227),
				.c(c2701K)
);

ninexnine_unit ninexnine_unit_5868(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2K008),
				.b1(W2K018),
				.b2(W2K028),
				.b3(W2K108),
				.b4(W2K118),
				.b5(W2K128),
				.b6(W2K208),
				.b7(W2K218),
				.b8(W2K228),
				.c(c2801K)
);

ninexnine_unit ninexnine_unit_5869(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2K009),
				.b1(W2K019),
				.b2(W2K029),
				.b3(W2K109),
				.b4(W2K119),
				.b5(W2K129),
				.b6(W2K209),
				.b7(W2K219),
				.b8(W2K229),
				.c(c2901K)
);

ninexnine_unit ninexnine_unit_5870(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2K00A),
				.b1(W2K01A),
				.b2(W2K02A),
				.b3(W2K10A),
				.b4(W2K11A),
				.b5(W2K12A),
				.b6(W2K20A),
				.b7(W2K21A),
				.b8(W2K22A),
				.c(c2A01K)
);

ninexnine_unit ninexnine_unit_5871(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2K00B),
				.b1(W2K01B),
				.b2(W2K02B),
				.b3(W2K10B),
				.b4(W2K11B),
				.b5(W2K12B),
				.b6(W2K20B),
				.b7(W2K21B),
				.b8(W2K22B),
				.c(c2B01K)
);

ninexnine_unit ninexnine_unit_5872(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2K00C),
				.b1(W2K01C),
				.b2(W2K02C),
				.b3(W2K10C),
				.b4(W2K11C),
				.b5(W2K12C),
				.b6(W2K20C),
				.b7(W2K21C),
				.b8(W2K22C),
				.c(c2C01K)
);

ninexnine_unit ninexnine_unit_5873(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2K00D),
				.b1(W2K01D),
				.b2(W2K02D),
				.b3(W2K10D),
				.b4(W2K11D),
				.b5(W2K12D),
				.b6(W2K20D),
				.b7(W2K21D),
				.b8(W2K22D),
				.c(c2D01K)
);

ninexnine_unit ninexnine_unit_5874(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2K00E),
				.b1(W2K01E),
				.b2(W2K02E),
				.b3(W2K10E),
				.b4(W2K11E),
				.b5(W2K12E),
				.b6(W2K20E),
				.b7(W2K21E),
				.b8(W2K22E),
				.c(c2E01K)
);

ninexnine_unit ninexnine_unit_5875(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2K00F),
				.b1(W2K01F),
				.b2(W2K02F),
				.b3(W2K10F),
				.b4(W2K11F),
				.b5(W2K12F),
				.b6(W2K20F),
				.b7(W2K21F),
				.b8(W2K22F),
				.c(c2F01K)
);

assign C201K=c2001K+c2101K+c2201K+c2301K+c2401K+c2501K+c2601K+c2701K+c2801K+c2901K+c2A01K+c2B01K+c2C01K+c2D01K+c2E01K+c2F01K;
assign A201K=(C201K>=0)?1:0;

assign P301K=A201K;

ninexnine_unit ninexnine_unit_5876(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2K000),
				.b1(W2K010),
				.b2(W2K020),
				.b3(W2K100),
				.b4(W2K110),
				.b5(W2K120),
				.b6(W2K200),
				.b7(W2K210),
				.b8(W2K220),
				.c(c2002K)
);

ninexnine_unit ninexnine_unit_5877(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2K001),
				.b1(W2K011),
				.b2(W2K021),
				.b3(W2K101),
				.b4(W2K111),
				.b5(W2K121),
				.b6(W2K201),
				.b7(W2K211),
				.b8(W2K221),
				.c(c2102K)
);

ninexnine_unit ninexnine_unit_5878(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2K002),
				.b1(W2K012),
				.b2(W2K022),
				.b3(W2K102),
				.b4(W2K112),
				.b5(W2K122),
				.b6(W2K202),
				.b7(W2K212),
				.b8(W2K222),
				.c(c2202K)
);

ninexnine_unit ninexnine_unit_5879(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2K003),
				.b1(W2K013),
				.b2(W2K023),
				.b3(W2K103),
				.b4(W2K113),
				.b5(W2K123),
				.b6(W2K203),
				.b7(W2K213),
				.b8(W2K223),
				.c(c2302K)
);

ninexnine_unit ninexnine_unit_5880(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2K004),
				.b1(W2K014),
				.b2(W2K024),
				.b3(W2K104),
				.b4(W2K114),
				.b5(W2K124),
				.b6(W2K204),
				.b7(W2K214),
				.b8(W2K224),
				.c(c2402K)
);

ninexnine_unit ninexnine_unit_5881(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2K005),
				.b1(W2K015),
				.b2(W2K025),
				.b3(W2K105),
				.b4(W2K115),
				.b5(W2K125),
				.b6(W2K205),
				.b7(W2K215),
				.b8(W2K225),
				.c(c2502K)
);

ninexnine_unit ninexnine_unit_5882(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2K006),
				.b1(W2K016),
				.b2(W2K026),
				.b3(W2K106),
				.b4(W2K116),
				.b5(W2K126),
				.b6(W2K206),
				.b7(W2K216),
				.b8(W2K226),
				.c(c2602K)
);

ninexnine_unit ninexnine_unit_5883(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2K007),
				.b1(W2K017),
				.b2(W2K027),
				.b3(W2K107),
				.b4(W2K117),
				.b5(W2K127),
				.b6(W2K207),
				.b7(W2K217),
				.b8(W2K227),
				.c(c2702K)
);

ninexnine_unit ninexnine_unit_5884(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2K008),
				.b1(W2K018),
				.b2(W2K028),
				.b3(W2K108),
				.b4(W2K118),
				.b5(W2K128),
				.b6(W2K208),
				.b7(W2K218),
				.b8(W2K228),
				.c(c2802K)
);

ninexnine_unit ninexnine_unit_5885(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2K009),
				.b1(W2K019),
				.b2(W2K029),
				.b3(W2K109),
				.b4(W2K119),
				.b5(W2K129),
				.b6(W2K209),
				.b7(W2K219),
				.b8(W2K229),
				.c(c2902K)
);

ninexnine_unit ninexnine_unit_5886(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2K00A),
				.b1(W2K01A),
				.b2(W2K02A),
				.b3(W2K10A),
				.b4(W2K11A),
				.b5(W2K12A),
				.b6(W2K20A),
				.b7(W2K21A),
				.b8(W2K22A),
				.c(c2A02K)
);

ninexnine_unit ninexnine_unit_5887(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2K00B),
				.b1(W2K01B),
				.b2(W2K02B),
				.b3(W2K10B),
				.b4(W2K11B),
				.b5(W2K12B),
				.b6(W2K20B),
				.b7(W2K21B),
				.b8(W2K22B),
				.c(c2B02K)
);

ninexnine_unit ninexnine_unit_5888(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2K00C),
				.b1(W2K01C),
				.b2(W2K02C),
				.b3(W2K10C),
				.b4(W2K11C),
				.b5(W2K12C),
				.b6(W2K20C),
				.b7(W2K21C),
				.b8(W2K22C),
				.c(c2C02K)
);

ninexnine_unit ninexnine_unit_5889(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2K00D),
				.b1(W2K01D),
				.b2(W2K02D),
				.b3(W2K10D),
				.b4(W2K11D),
				.b5(W2K12D),
				.b6(W2K20D),
				.b7(W2K21D),
				.b8(W2K22D),
				.c(c2D02K)
);

ninexnine_unit ninexnine_unit_5890(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2K00E),
				.b1(W2K01E),
				.b2(W2K02E),
				.b3(W2K10E),
				.b4(W2K11E),
				.b5(W2K12E),
				.b6(W2K20E),
				.b7(W2K21E),
				.b8(W2K22E),
				.c(c2E02K)
);

ninexnine_unit ninexnine_unit_5891(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2K00F),
				.b1(W2K01F),
				.b2(W2K02F),
				.b3(W2K10F),
				.b4(W2K11F),
				.b5(W2K12F),
				.b6(W2K20F),
				.b7(W2K21F),
				.b8(W2K22F),
				.c(c2F02K)
);

assign C202K=c2002K+c2102K+c2202K+c2302K+c2402K+c2502K+c2602K+c2702K+c2802K+c2902K+c2A02K+c2B02K+c2C02K+c2D02K+c2E02K+c2F02K;
assign A202K=(C202K>=0)?1:0;

assign P302K=A202K;

ninexnine_unit ninexnine_unit_5892(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2K000),
				.b1(W2K010),
				.b2(W2K020),
				.b3(W2K100),
				.b4(W2K110),
				.b5(W2K120),
				.b6(W2K200),
				.b7(W2K210),
				.b8(W2K220),
				.c(c2010K)
);

ninexnine_unit ninexnine_unit_5893(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2K001),
				.b1(W2K011),
				.b2(W2K021),
				.b3(W2K101),
				.b4(W2K111),
				.b5(W2K121),
				.b6(W2K201),
				.b7(W2K211),
				.b8(W2K221),
				.c(c2110K)
);

ninexnine_unit ninexnine_unit_5894(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2K002),
				.b1(W2K012),
				.b2(W2K022),
				.b3(W2K102),
				.b4(W2K112),
				.b5(W2K122),
				.b6(W2K202),
				.b7(W2K212),
				.b8(W2K222),
				.c(c2210K)
);

ninexnine_unit ninexnine_unit_5895(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2K003),
				.b1(W2K013),
				.b2(W2K023),
				.b3(W2K103),
				.b4(W2K113),
				.b5(W2K123),
				.b6(W2K203),
				.b7(W2K213),
				.b8(W2K223),
				.c(c2310K)
);

ninexnine_unit ninexnine_unit_5896(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2K004),
				.b1(W2K014),
				.b2(W2K024),
				.b3(W2K104),
				.b4(W2K114),
				.b5(W2K124),
				.b6(W2K204),
				.b7(W2K214),
				.b8(W2K224),
				.c(c2410K)
);

ninexnine_unit ninexnine_unit_5897(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2K005),
				.b1(W2K015),
				.b2(W2K025),
				.b3(W2K105),
				.b4(W2K115),
				.b5(W2K125),
				.b6(W2K205),
				.b7(W2K215),
				.b8(W2K225),
				.c(c2510K)
);

ninexnine_unit ninexnine_unit_5898(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2K006),
				.b1(W2K016),
				.b2(W2K026),
				.b3(W2K106),
				.b4(W2K116),
				.b5(W2K126),
				.b6(W2K206),
				.b7(W2K216),
				.b8(W2K226),
				.c(c2610K)
);

ninexnine_unit ninexnine_unit_5899(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2K007),
				.b1(W2K017),
				.b2(W2K027),
				.b3(W2K107),
				.b4(W2K117),
				.b5(W2K127),
				.b6(W2K207),
				.b7(W2K217),
				.b8(W2K227),
				.c(c2710K)
);

ninexnine_unit ninexnine_unit_5900(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2K008),
				.b1(W2K018),
				.b2(W2K028),
				.b3(W2K108),
				.b4(W2K118),
				.b5(W2K128),
				.b6(W2K208),
				.b7(W2K218),
				.b8(W2K228),
				.c(c2810K)
);

ninexnine_unit ninexnine_unit_5901(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2K009),
				.b1(W2K019),
				.b2(W2K029),
				.b3(W2K109),
				.b4(W2K119),
				.b5(W2K129),
				.b6(W2K209),
				.b7(W2K219),
				.b8(W2K229),
				.c(c2910K)
);

ninexnine_unit ninexnine_unit_5902(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2K00A),
				.b1(W2K01A),
				.b2(W2K02A),
				.b3(W2K10A),
				.b4(W2K11A),
				.b5(W2K12A),
				.b6(W2K20A),
				.b7(W2K21A),
				.b8(W2K22A),
				.c(c2A10K)
);

ninexnine_unit ninexnine_unit_5903(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2K00B),
				.b1(W2K01B),
				.b2(W2K02B),
				.b3(W2K10B),
				.b4(W2K11B),
				.b5(W2K12B),
				.b6(W2K20B),
				.b7(W2K21B),
				.b8(W2K22B),
				.c(c2B10K)
);

ninexnine_unit ninexnine_unit_5904(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2K00C),
				.b1(W2K01C),
				.b2(W2K02C),
				.b3(W2K10C),
				.b4(W2K11C),
				.b5(W2K12C),
				.b6(W2K20C),
				.b7(W2K21C),
				.b8(W2K22C),
				.c(c2C10K)
);

ninexnine_unit ninexnine_unit_5905(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2K00D),
				.b1(W2K01D),
				.b2(W2K02D),
				.b3(W2K10D),
				.b4(W2K11D),
				.b5(W2K12D),
				.b6(W2K20D),
				.b7(W2K21D),
				.b8(W2K22D),
				.c(c2D10K)
);

ninexnine_unit ninexnine_unit_5906(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2K00E),
				.b1(W2K01E),
				.b2(W2K02E),
				.b3(W2K10E),
				.b4(W2K11E),
				.b5(W2K12E),
				.b6(W2K20E),
				.b7(W2K21E),
				.b8(W2K22E),
				.c(c2E10K)
);

ninexnine_unit ninexnine_unit_5907(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2K00F),
				.b1(W2K01F),
				.b2(W2K02F),
				.b3(W2K10F),
				.b4(W2K11F),
				.b5(W2K12F),
				.b6(W2K20F),
				.b7(W2K21F),
				.b8(W2K22F),
				.c(c2F10K)
);

assign C210K=c2010K+c2110K+c2210K+c2310K+c2410K+c2510K+c2610K+c2710K+c2810K+c2910K+c2A10K+c2B10K+c2C10K+c2D10K+c2E10K+c2F10K;
assign A210K=(C210K>=0)?1:0;

assign P310K=A210K;

ninexnine_unit ninexnine_unit_5908(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2K000),
				.b1(W2K010),
				.b2(W2K020),
				.b3(W2K100),
				.b4(W2K110),
				.b5(W2K120),
				.b6(W2K200),
				.b7(W2K210),
				.b8(W2K220),
				.c(c2011K)
);

ninexnine_unit ninexnine_unit_5909(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2K001),
				.b1(W2K011),
				.b2(W2K021),
				.b3(W2K101),
				.b4(W2K111),
				.b5(W2K121),
				.b6(W2K201),
				.b7(W2K211),
				.b8(W2K221),
				.c(c2111K)
);

ninexnine_unit ninexnine_unit_5910(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2K002),
				.b1(W2K012),
				.b2(W2K022),
				.b3(W2K102),
				.b4(W2K112),
				.b5(W2K122),
				.b6(W2K202),
				.b7(W2K212),
				.b8(W2K222),
				.c(c2211K)
);

ninexnine_unit ninexnine_unit_5911(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2K003),
				.b1(W2K013),
				.b2(W2K023),
				.b3(W2K103),
				.b4(W2K113),
				.b5(W2K123),
				.b6(W2K203),
				.b7(W2K213),
				.b8(W2K223),
				.c(c2311K)
);

ninexnine_unit ninexnine_unit_5912(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2K004),
				.b1(W2K014),
				.b2(W2K024),
				.b3(W2K104),
				.b4(W2K114),
				.b5(W2K124),
				.b6(W2K204),
				.b7(W2K214),
				.b8(W2K224),
				.c(c2411K)
);

ninexnine_unit ninexnine_unit_5913(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2K005),
				.b1(W2K015),
				.b2(W2K025),
				.b3(W2K105),
				.b4(W2K115),
				.b5(W2K125),
				.b6(W2K205),
				.b7(W2K215),
				.b8(W2K225),
				.c(c2511K)
);

ninexnine_unit ninexnine_unit_5914(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2K006),
				.b1(W2K016),
				.b2(W2K026),
				.b3(W2K106),
				.b4(W2K116),
				.b5(W2K126),
				.b6(W2K206),
				.b7(W2K216),
				.b8(W2K226),
				.c(c2611K)
);

ninexnine_unit ninexnine_unit_5915(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2K007),
				.b1(W2K017),
				.b2(W2K027),
				.b3(W2K107),
				.b4(W2K117),
				.b5(W2K127),
				.b6(W2K207),
				.b7(W2K217),
				.b8(W2K227),
				.c(c2711K)
);

ninexnine_unit ninexnine_unit_5916(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2K008),
				.b1(W2K018),
				.b2(W2K028),
				.b3(W2K108),
				.b4(W2K118),
				.b5(W2K128),
				.b6(W2K208),
				.b7(W2K218),
				.b8(W2K228),
				.c(c2811K)
);

ninexnine_unit ninexnine_unit_5917(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2K009),
				.b1(W2K019),
				.b2(W2K029),
				.b3(W2K109),
				.b4(W2K119),
				.b5(W2K129),
				.b6(W2K209),
				.b7(W2K219),
				.b8(W2K229),
				.c(c2911K)
);

ninexnine_unit ninexnine_unit_5918(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2K00A),
				.b1(W2K01A),
				.b2(W2K02A),
				.b3(W2K10A),
				.b4(W2K11A),
				.b5(W2K12A),
				.b6(W2K20A),
				.b7(W2K21A),
				.b8(W2K22A),
				.c(c2A11K)
);

ninexnine_unit ninexnine_unit_5919(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2K00B),
				.b1(W2K01B),
				.b2(W2K02B),
				.b3(W2K10B),
				.b4(W2K11B),
				.b5(W2K12B),
				.b6(W2K20B),
				.b7(W2K21B),
				.b8(W2K22B),
				.c(c2B11K)
);

ninexnine_unit ninexnine_unit_5920(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2K00C),
				.b1(W2K01C),
				.b2(W2K02C),
				.b3(W2K10C),
				.b4(W2K11C),
				.b5(W2K12C),
				.b6(W2K20C),
				.b7(W2K21C),
				.b8(W2K22C),
				.c(c2C11K)
);

ninexnine_unit ninexnine_unit_5921(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2K00D),
				.b1(W2K01D),
				.b2(W2K02D),
				.b3(W2K10D),
				.b4(W2K11D),
				.b5(W2K12D),
				.b6(W2K20D),
				.b7(W2K21D),
				.b8(W2K22D),
				.c(c2D11K)
);

ninexnine_unit ninexnine_unit_5922(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2K00E),
				.b1(W2K01E),
				.b2(W2K02E),
				.b3(W2K10E),
				.b4(W2K11E),
				.b5(W2K12E),
				.b6(W2K20E),
				.b7(W2K21E),
				.b8(W2K22E),
				.c(c2E11K)
);

ninexnine_unit ninexnine_unit_5923(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2K00F),
				.b1(W2K01F),
				.b2(W2K02F),
				.b3(W2K10F),
				.b4(W2K11F),
				.b5(W2K12F),
				.b6(W2K20F),
				.b7(W2K21F),
				.b8(W2K22F),
				.c(c2F11K)
);

assign C211K=c2011K+c2111K+c2211K+c2311K+c2411K+c2511K+c2611K+c2711K+c2811K+c2911K+c2A11K+c2B11K+c2C11K+c2D11K+c2E11K+c2F11K;
assign A211K=(C211K>=0)?1:0;

assign P311K=A211K;

ninexnine_unit ninexnine_unit_5924(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2K000),
				.b1(W2K010),
				.b2(W2K020),
				.b3(W2K100),
				.b4(W2K110),
				.b5(W2K120),
				.b6(W2K200),
				.b7(W2K210),
				.b8(W2K220),
				.c(c2012K)
);

ninexnine_unit ninexnine_unit_5925(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2K001),
				.b1(W2K011),
				.b2(W2K021),
				.b3(W2K101),
				.b4(W2K111),
				.b5(W2K121),
				.b6(W2K201),
				.b7(W2K211),
				.b8(W2K221),
				.c(c2112K)
);

ninexnine_unit ninexnine_unit_5926(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2K002),
				.b1(W2K012),
				.b2(W2K022),
				.b3(W2K102),
				.b4(W2K112),
				.b5(W2K122),
				.b6(W2K202),
				.b7(W2K212),
				.b8(W2K222),
				.c(c2212K)
);

ninexnine_unit ninexnine_unit_5927(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2K003),
				.b1(W2K013),
				.b2(W2K023),
				.b3(W2K103),
				.b4(W2K113),
				.b5(W2K123),
				.b6(W2K203),
				.b7(W2K213),
				.b8(W2K223),
				.c(c2312K)
);

ninexnine_unit ninexnine_unit_5928(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2K004),
				.b1(W2K014),
				.b2(W2K024),
				.b3(W2K104),
				.b4(W2K114),
				.b5(W2K124),
				.b6(W2K204),
				.b7(W2K214),
				.b8(W2K224),
				.c(c2412K)
);

ninexnine_unit ninexnine_unit_5929(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2K005),
				.b1(W2K015),
				.b2(W2K025),
				.b3(W2K105),
				.b4(W2K115),
				.b5(W2K125),
				.b6(W2K205),
				.b7(W2K215),
				.b8(W2K225),
				.c(c2512K)
);

ninexnine_unit ninexnine_unit_5930(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2K006),
				.b1(W2K016),
				.b2(W2K026),
				.b3(W2K106),
				.b4(W2K116),
				.b5(W2K126),
				.b6(W2K206),
				.b7(W2K216),
				.b8(W2K226),
				.c(c2612K)
);

ninexnine_unit ninexnine_unit_5931(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2K007),
				.b1(W2K017),
				.b2(W2K027),
				.b3(W2K107),
				.b4(W2K117),
				.b5(W2K127),
				.b6(W2K207),
				.b7(W2K217),
				.b8(W2K227),
				.c(c2712K)
);

ninexnine_unit ninexnine_unit_5932(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2K008),
				.b1(W2K018),
				.b2(W2K028),
				.b3(W2K108),
				.b4(W2K118),
				.b5(W2K128),
				.b6(W2K208),
				.b7(W2K218),
				.b8(W2K228),
				.c(c2812K)
);

ninexnine_unit ninexnine_unit_5933(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2K009),
				.b1(W2K019),
				.b2(W2K029),
				.b3(W2K109),
				.b4(W2K119),
				.b5(W2K129),
				.b6(W2K209),
				.b7(W2K219),
				.b8(W2K229),
				.c(c2912K)
);

ninexnine_unit ninexnine_unit_5934(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2K00A),
				.b1(W2K01A),
				.b2(W2K02A),
				.b3(W2K10A),
				.b4(W2K11A),
				.b5(W2K12A),
				.b6(W2K20A),
				.b7(W2K21A),
				.b8(W2K22A),
				.c(c2A12K)
);

ninexnine_unit ninexnine_unit_5935(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2K00B),
				.b1(W2K01B),
				.b2(W2K02B),
				.b3(W2K10B),
				.b4(W2K11B),
				.b5(W2K12B),
				.b6(W2K20B),
				.b7(W2K21B),
				.b8(W2K22B),
				.c(c2B12K)
);

ninexnine_unit ninexnine_unit_5936(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2K00C),
				.b1(W2K01C),
				.b2(W2K02C),
				.b3(W2K10C),
				.b4(W2K11C),
				.b5(W2K12C),
				.b6(W2K20C),
				.b7(W2K21C),
				.b8(W2K22C),
				.c(c2C12K)
);

ninexnine_unit ninexnine_unit_5937(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2K00D),
				.b1(W2K01D),
				.b2(W2K02D),
				.b3(W2K10D),
				.b4(W2K11D),
				.b5(W2K12D),
				.b6(W2K20D),
				.b7(W2K21D),
				.b8(W2K22D),
				.c(c2D12K)
);

ninexnine_unit ninexnine_unit_5938(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2K00E),
				.b1(W2K01E),
				.b2(W2K02E),
				.b3(W2K10E),
				.b4(W2K11E),
				.b5(W2K12E),
				.b6(W2K20E),
				.b7(W2K21E),
				.b8(W2K22E),
				.c(c2E12K)
);

ninexnine_unit ninexnine_unit_5939(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2K00F),
				.b1(W2K01F),
				.b2(W2K02F),
				.b3(W2K10F),
				.b4(W2K11F),
				.b5(W2K12F),
				.b6(W2K20F),
				.b7(W2K21F),
				.b8(W2K22F),
				.c(c2F12K)
);

assign C212K=c2012K+c2112K+c2212K+c2312K+c2412K+c2512K+c2612K+c2712K+c2812K+c2912K+c2A12K+c2B12K+c2C12K+c2D12K+c2E12K+c2F12K;
assign A212K=(C212K>=0)?1:0;

assign P312K=A212K;

ninexnine_unit ninexnine_unit_5940(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2K000),
				.b1(W2K010),
				.b2(W2K020),
				.b3(W2K100),
				.b4(W2K110),
				.b5(W2K120),
				.b6(W2K200),
				.b7(W2K210),
				.b8(W2K220),
				.c(c2020K)
);

ninexnine_unit ninexnine_unit_5941(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2K001),
				.b1(W2K011),
				.b2(W2K021),
				.b3(W2K101),
				.b4(W2K111),
				.b5(W2K121),
				.b6(W2K201),
				.b7(W2K211),
				.b8(W2K221),
				.c(c2120K)
);

ninexnine_unit ninexnine_unit_5942(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2K002),
				.b1(W2K012),
				.b2(W2K022),
				.b3(W2K102),
				.b4(W2K112),
				.b5(W2K122),
				.b6(W2K202),
				.b7(W2K212),
				.b8(W2K222),
				.c(c2220K)
);

ninexnine_unit ninexnine_unit_5943(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2K003),
				.b1(W2K013),
				.b2(W2K023),
				.b3(W2K103),
				.b4(W2K113),
				.b5(W2K123),
				.b6(W2K203),
				.b7(W2K213),
				.b8(W2K223),
				.c(c2320K)
);

ninexnine_unit ninexnine_unit_5944(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2K004),
				.b1(W2K014),
				.b2(W2K024),
				.b3(W2K104),
				.b4(W2K114),
				.b5(W2K124),
				.b6(W2K204),
				.b7(W2K214),
				.b8(W2K224),
				.c(c2420K)
);

ninexnine_unit ninexnine_unit_5945(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2K005),
				.b1(W2K015),
				.b2(W2K025),
				.b3(W2K105),
				.b4(W2K115),
				.b5(W2K125),
				.b6(W2K205),
				.b7(W2K215),
				.b8(W2K225),
				.c(c2520K)
);

ninexnine_unit ninexnine_unit_5946(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2K006),
				.b1(W2K016),
				.b2(W2K026),
				.b3(W2K106),
				.b4(W2K116),
				.b5(W2K126),
				.b6(W2K206),
				.b7(W2K216),
				.b8(W2K226),
				.c(c2620K)
);

ninexnine_unit ninexnine_unit_5947(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2K007),
				.b1(W2K017),
				.b2(W2K027),
				.b3(W2K107),
				.b4(W2K117),
				.b5(W2K127),
				.b6(W2K207),
				.b7(W2K217),
				.b8(W2K227),
				.c(c2720K)
);

ninexnine_unit ninexnine_unit_5948(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2K008),
				.b1(W2K018),
				.b2(W2K028),
				.b3(W2K108),
				.b4(W2K118),
				.b5(W2K128),
				.b6(W2K208),
				.b7(W2K218),
				.b8(W2K228),
				.c(c2820K)
);

ninexnine_unit ninexnine_unit_5949(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2K009),
				.b1(W2K019),
				.b2(W2K029),
				.b3(W2K109),
				.b4(W2K119),
				.b5(W2K129),
				.b6(W2K209),
				.b7(W2K219),
				.b8(W2K229),
				.c(c2920K)
);

ninexnine_unit ninexnine_unit_5950(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2K00A),
				.b1(W2K01A),
				.b2(W2K02A),
				.b3(W2K10A),
				.b4(W2K11A),
				.b5(W2K12A),
				.b6(W2K20A),
				.b7(W2K21A),
				.b8(W2K22A),
				.c(c2A20K)
);

ninexnine_unit ninexnine_unit_5951(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2K00B),
				.b1(W2K01B),
				.b2(W2K02B),
				.b3(W2K10B),
				.b4(W2K11B),
				.b5(W2K12B),
				.b6(W2K20B),
				.b7(W2K21B),
				.b8(W2K22B),
				.c(c2B20K)
);

ninexnine_unit ninexnine_unit_5952(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2K00C),
				.b1(W2K01C),
				.b2(W2K02C),
				.b3(W2K10C),
				.b4(W2K11C),
				.b5(W2K12C),
				.b6(W2K20C),
				.b7(W2K21C),
				.b8(W2K22C),
				.c(c2C20K)
);

ninexnine_unit ninexnine_unit_5953(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2K00D),
				.b1(W2K01D),
				.b2(W2K02D),
				.b3(W2K10D),
				.b4(W2K11D),
				.b5(W2K12D),
				.b6(W2K20D),
				.b7(W2K21D),
				.b8(W2K22D),
				.c(c2D20K)
);

ninexnine_unit ninexnine_unit_5954(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2K00E),
				.b1(W2K01E),
				.b2(W2K02E),
				.b3(W2K10E),
				.b4(W2K11E),
				.b5(W2K12E),
				.b6(W2K20E),
				.b7(W2K21E),
				.b8(W2K22E),
				.c(c2E20K)
);

ninexnine_unit ninexnine_unit_5955(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2K00F),
				.b1(W2K01F),
				.b2(W2K02F),
				.b3(W2K10F),
				.b4(W2K11F),
				.b5(W2K12F),
				.b6(W2K20F),
				.b7(W2K21F),
				.b8(W2K22F),
				.c(c2F20K)
);

assign C220K=c2020K+c2120K+c2220K+c2320K+c2420K+c2520K+c2620K+c2720K+c2820K+c2920K+c2A20K+c2B20K+c2C20K+c2D20K+c2E20K+c2F20K;
assign A220K=(C220K>=0)?1:0;

assign P320K=A220K;

ninexnine_unit ninexnine_unit_5956(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2K000),
				.b1(W2K010),
				.b2(W2K020),
				.b3(W2K100),
				.b4(W2K110),
				.b5(W2K120),
				.b6(W2K200),
				.b7(W2K210),
				.b8(W2K220),
				.c(c2021K)
);

ninexnine_unit ninexnine_unit_5957(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2K001),
				.b1(W2K011),
				.b2(W2K021),
				.b3(W2K101),
				.b4(W2K111),
				.b5(W2K121),
				.b6(W2K201),
				.b7(W2K211),
				.b8(W2K221),
				.c(c2121K)
);

ninexnine_unit ninexnine_unit_5958(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2K002),
				.b1(W2K012),
				.b2(W2K022),
				.b3(W2K102),
				.b4(W2K112),
				.b5(W2K122),
				.b6(W2K202),
				.b7(W2K212),
				.b8(W2K222),
				.c(c2221K)
);

ninexnine_unit ninexnine_unit_5959(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2K003),
				.b1(W2K013),
				.b2(W2K023),
				.b3(W2K103),
				.b4(W2K113),
				.b5(W2K123),
				.b6(W2K203),
				.b7(W2K213),
				.b8(W2K223),
				.c(c2321K)
);

ninexnine_unit ninexnine_unit_5960(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2K004),
				.b1(W2K014),
				.b2(W2K024),
				.b3(W2K104),
				.b4(W2K114),
				.b5(W2K124),
				.b6(W2K204),
				.b7(W2K214),
				.b8(W2K224),
				.c(c2421K)
);

ninexnine_unit ninexnine_unit_5961(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2K005),
				.b1(W2K015),
				.b2(W2K025),
				.b3(W2K105),
				.b4(W2K115),
				.b5(W2K125),
				.b6(W2K205),
				.b7(W2K215),
				.b8(W2K225),
				.c(c2521K)
);

ninexnine_unit ninexnine_unit_5962(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2K006),
				.b1(W2K016),
				.b2(W2K026),
				.b3(W2K106),
				.b4(W2K116),
				.b5(W2K126),
				.b6(W2K206),
				.b7(W2K216),
				.b8(W2K226),
				.c(c2621K)
);

ninexnine_unit ninexnine_unit_5963(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2K007),
				.b1(W2K017),
				.b2(W2K027),
				.b3(W2K107),
				.b4(W2K117),
				.b5(W2K127),
				.b6(W2K207),
				.b7(W2K217),
				.b8(W2K227),
				.c(c2721K)
);

ninexnine_unit ninexnine_unit_5964(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2K008),
				.b1(W2K018),
				.b2(W2K028),
				.b3(W2K108),
				.b4(W2K118),
				.b5(W2K128),
				.b6(W2K208),
				.b7(W2K218),
				.b8(W2K228),
				.c(c2821K)
);

ninexnine_unit ninexnine_unit_5965(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2K009),
				.b1(W2K019),
				.b2(W2K029),
				.b3(W2K109),
				.b4(W2K119),
				.b5(W2K129),
				.b6(W2K209),
				.b7(W2K219),
				.b8(W2K229),
				.c(c2921K)
);

ninexnine_unit ninexnine_unit_5966(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2K00A),
				.b1(W2K01A),
				.b2(W2K02A),
				.b3(W2K10A),
				.b4(W2K11A),
				.b5(W2K12A),
				.b6(W2K20A),
				.b7(W2K21A),
				.b8(W2K22A),
				.c(c2A21K)
);

ninexnine_unit ninexnine_unit_5967(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2K00B),
				.b1(W2K01B),
				.b2(W2K02B),
				.b3(W2K10B),
				.b4(W2K11B),
				.b5(W2K12B),
				.b6(W2K20B),
				.b7(W2K21B),
				.b8(W2K22B),
				.c(c2B21K)
);

ninexnine_unit ninexnine_unit_5968(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2K00C),
				.b1(W2K01C),
				.b2(W2K02C),
				.b3(W2K10C),
				.b4(W2K11C),
				.b5(W2K12C),
				.b6(W2K20C),
				.b7(W2K21C),
				.b8(W2K22C),
				.c(c2C21K)
);

ninexnine_unit ninexnine_unit_5969(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2K00D),
				.b1(W2K01D),
				.b2(W2K02D),
				.b3(W2K10D),
				.b4(W2K11D),
				.b5(W2K12D),
				.b6(W2K20D),
				.b7(W2K21D),
				.b8(W2K22D),
				.c(c2D21K)
);

ninexnine_unit ninexnine_unit_5970(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2K00E),
				.b1(W2K01E),
				.b2(W2K02E),
				.b3(W2K10E),
				.b4(W2K11E),
				.b5(W2K12E),
				.b6(W2K20E),
				.b7(W2K21E),
				.b8(W2K22E),
				.c(c2E21K)
);

ninexnine_unit ninexnine_unit_5971(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2K00F),
				.b1(W2K01F),
				.b2(W2K02F),
				.b3(W2K10F),
				.b4(W2K11F),
				.b5(W2K12F),
				.b6(W2K20F),
				.b7(W2K21F),
				.b8(W2K22F),
				.c(c2F21K)
);

assign C221K=c2021K+c2121K+c2221K+c2321K+c2421K+c2521K+c2621K+c2721K+c2821K+c2921K+c2A21K+c2B21K+c2C21K+c2D21K+c2E21K+c2F21K;
assign A221K=(C221K>=0)?1:0;

assign P321K=A221K;

ninexnine_unit ninexnine_unit_5972(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2K000),
				.b1(W2K010),
				.b2(W2K020),
				.b3(W2K100),
				.b4(W2K110),
				.b5(W2K120),
				.b6(W2K200),
				.b7(W2K210),
				.b8(W2K220),
				.c(c2022K)
);

ninexnine_unit ninexnine_unit_5973(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2K001),
				.b1(W2K011),
				.b2(W2K021),
				.b3(W2K101),
				.b4(W2K111),
				.b5(W2K121),
				.b6(W2K201),
				.b7(W2K211),
				.b8(W2K221),
				.c(c2122K)
);

ninexnine_unit ninexnine_unit_5974(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2K002),
				.b1(W2K012),
				.b2(W2K022),
				.b3(W2K102),
				.b4(W2K112),
				.b5(W2K122),
				.b6(W2K202),
				.b7(W2K212),
				.b8(W2K222),
				.c(c2222K)
);

ninexnine_unit ninexnine_unit_5975(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2K003),
				.b1(W2K013),
				.b2(W2K023),
				.b3(W2K103),
				.b4(W2K113),
				.b5(W2K123),
				.b6(W2K203),
				.b7(W2K213),
				.b8(W2K223),
				.c(c2322K)
);

ninexnine_unit ninexnine_unit_5976(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2K004),
				.b1(W2K014),
				.b2(W2K024),
				.b3(W2K104),
				.b4(W2K114),
				.b5(W2K124),
				.b6(W2K204),
				.b7(W2K214),
				.b8(W2K224),
				.c(c2422K)
);

ninexnine_unit ninexnine_unit_5977(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2K005),
				.b1(W2K015),
				.b2(W2K025),
				.b3(W2K105),
				.b4(W2K115),
				.b5(W2K125),
				.b6(W2K205),
				.b7(W2K215),
				.b8(W2K225),
				.c(c2522K)
);

ninexnine_unit ninexnine_unit_5978(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2K006),
				.b1(W2K016),
				.b2(W2K026),
				.b3(W2K106),
				.b4(W2K116),
				.b5(W2K126),
				.b6(W2K206),
				.b7(W2K216),
				.b8(W2K226),
				.c(c2622K)
);

ninexnine_unit ninexnine_unit_5979(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2K007),
				.b1(W2K017),
				.b2(W2K027),
				.b3(W2K107),
				.b4(W2K117),
				.b5(W2K127),
				.b6(W2K207),
				.b7(W2K217),
				.b8(W2K227),
				.c(c2722K)
);

ninexnine_unit ninexnine_unit_5980(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2K008),
				.b1(W2K018),
				.b2(W2K028),
				.b3(W2K108),
				.b4(W2K118),
				.b5(W2K128),
				.b6(W2K208),
				.b7(W2K218),
				.b8(W2K228),
				.c(c2822K)
);

ninexnine_unit ninexnine_unit_5981(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2K009),
				.b1(W2K019),
				.b2(W2K029),
				.b3(W2K109),
				.b4(W2K119),
				.b5(W2K129),
				.b6(W2K209),
				.b7(W2K219),
				.b8(W2K229),
				.c(c2922K)
);

ninexnine_unit ninexnine_unit_5982(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2K00A),
				.b1(W2K01A),
				.b2(W2K02A),
				.b3(W2K10A),
				.b4(W2K11A),
				.b5(W2K12A),
				.b6(W2K20A),
				.b7(W2K21A),
				.b8(W2K22A),
				.c(c2A22K)
);

ninexnine_unit ninexnine_unit_5983(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2K00B),
				.b1(W2K01B),
				.b2(W2K02B),
				.b3(W2K10B),
				.b4(W2K11B),
				.b5(W2K12B),
				.b6(W2K20B),
				.b7(W2K21B),
				.b8(W2K22B),
				.c(c2B22K)
);

ninexnine_unit ninexnine_unit_5984(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2K00C),
				.b1(W2K01C),
				.b2(W2K02C),
				.b3(W2K10C),
				.b4(W2K11C),
				.b5(W2K12C),
				.b6(W2K20C),
				.b7(W2K21C),
				.b8(W2K22C),
				.c(c2C22K)
);

ninexnine_unit ninexnine_unit_5985(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2K00D),
				.b1(W2K01D),
				.b2(W2K02D),
				.b3(W2K10D),
				.b4(W2K11D),
				.b5(W2K12D),
				.b6(W2K20D),
				.b7(W2K21D),
				.b8(W2K22D),
				.c(c2D22K)
);

ninexnine_unit ninexnine_unit_5986(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2K00E),
				.b1(W2K01E),
				.b2(W2K02E),
				.b3(W2K10E),
				.b4(W2K11E),
				.b5(W2K12E),
				.b6(W2K20E),
				.b7(W2K21E),
				.b8(W2K22E),
				.c(c2E22K)
);

ninexnine_unit ninexnine_unit_5987(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2K00F),
				.b1(W2K01F),
				.b2(W2K02F),
				.b3(W2K10F),
				.b4(W2K11F),
				.b5(W2K12F),
				.b6(W2K20F),
				.b7(W2K21F),
				.b8(W2K22F),
				.c(c2F22K)
);

assign C222K=c2022K+c2122K+c2222K+c2322K+c2422K+c2522K+c2622K+c2722K+c2822K+c2922K+c2A22K+c2B22K+c2C22K+c2D22K+c2E22K+c2F22K;
assign A222K=(C222K>=0)?1:0;

assign P322K=A222K;

ninexnine_unit ninexnine_unit_5988(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2L000),
				.b1(W2L010),
				.b2(W2L020),
				.b3(W2L100),
				.b4(W2L110),
				.b5(W2L120),
				.b6(W2L200),
				.b7(W2L210),
				.b8(W2L220),
				.c(c2000L)
);

ninexnine_unit ninexnine_unit_5989(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2L001),
				.b1(W2L011),
				.b2(W2L021),
				.b3(W2L101),
				.b4(W2L111),
				.b5(W2L121),
				.b6(W2L201),
				.b7(W2L211),
				.b8(W2L221),
				.c(c2100L)
);

ninexnine_unit ninexnine_unit_5990(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2L002),
				.b1(W2L012),
				.b2(W2L022),
				.b3(W2L102),
				.b4(W2L112),
				.b5(W2L122),
				.b6(W2L202),
				.b7(W2L212),
				.b8(W2L222),
				.c(c2200L)
);

ninexnine_unit ninexnine_unit_5991(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2L003),
				.b1(W2L013),
				.b2(W2L023),
				.b3(W2L103),
				.b4(W2L113),
				.b5(W2L123),
				.b6(W2L203),
				.b7(W2L213),
				.b8(W2L223),
				.c(c2300L)
);

ninexnine_unit ninexnine_unit_5992(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2L004),
				.b1(W2L014),
				.b2(W2L024),
				.b3(W2L104),
				.b4(W2L114),
				.b5(W2L124),
				.b6(W2L204),
				.b7(W2L214),
				.b8(W2L224),
				.c(c2400L)
);

ninexnine_unit ninexnine_unit_5993(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2L005),
				.b1(W2L015),
				.b2(W2L025),
				.b3(W2L105),
				.b4(W2L115),
				.b5(W2L125),
				.b6(W2L205),
				.b7(W2L215),
				.b8(W2L225),
				.c(c2500L)
);

ninexnine_unit ninexnine_unit_5994(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2L006),
				.b1(W2L016),
				.b2(W2L026),
				.b3(W2L106),
				.b4(W2L116),
				.b5(W2L126),
				.b6(W2L206),
				.b7(W2L216),
				.b8(W2L226),
				.c(c2600L)
);

ninexnine_unit ninexnine_unit_5995(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2L007),
				.b1(W2L017),
				.b2(W2L027),
				.b3(W2L107),
				.b4(W2L117),
				.b5(W2L127),
				.b6(W2L207),
				.b7(W2L217),
				.b8(W2L227),
				.c(c2700L)
);

ninexnine_unit ninexnine_unit_5996(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2L008),
				.b1(W2L018),
				.b2(W2L028),
				.b3(W2L108),
				.b4(W2L118),
				.b5(W2L128),
				.b6(W2L208),
				.b7(W2L218),
				.b8(W2L228),
				.c(c2800L)
);

ninexnine_unit ninexnine_unit_5997(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2L009),
				.b1(W2L019),
				.b2(W2L029),
				.b3(W2L109),
				.b4(W2L119),
				.b5(W2L129),
				.b6(W2L209),
				.b7(W2L219),
				.b8(W2L229),
				.c(c2900L)
);

ninexnine_unit ninexnine_unit_5998(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2L00A),
				.b1(W2L01A),
				.b2(W2L02A),
				.b3(W2L10A),
				.b4(W2L11A),
				.b5(W2L12A),
				.b6(W2L20A),
				.b7(W2L21A),
				.b8(W2L22A),
				.c(c2A00L)
);

ninexnine_unit ninexnine_unit_5999(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2L00B),
				.b1(W2L01B),
				.b2(W2L02B),
				.b3(W2L10B),
				.b4(W2L11B),
				.b5(W2L12B),
				.b6(W2L20B),
				.b7(W2L21B),
				.b8(W2L22B),
				.c(c2B00L)
);

ninexnine_unit ninexnine_unit_6000(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2L00C),
				.b1(W2L01C),
				.b2(W2L02C),
				.b3(W2L10C),
				.b4(W2L11C),
				.b5(W2L12C),
				.b6(W2L20C),
				.b7(W2L21C),
				.b8(W2L22C),
				.c(c2C00L)
);

ninexnine_unit ninexnine_unit_6001(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2L00D),
				.b1(W2L01D),
				.b2(W2L02D),
				.b3(W2L10D),
				.b4(W2L11D),
				.b5(W2L12D),
				.b6(W2L20D),
				.b7(W2L21D),
				.b8(W2L22D),
				.c(c2D00L)
);

ninexnine_unit ninexnine_unit_6002(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2L00E),
				.b1(W2L01E),
				.b2(W2L02E),
				.b3(W2L10E),
				.b4(W2L11E),
				.b5(W2L12E),
				.b6(W2L20E),
				.b7(W2L21E),
				.b8(W2L22E),
				.c(c2E00L)
);

ninexnine_unit ninexnine_unit_6003(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2L00F),
				.b1(W2L01F),
				.b2(W2L02F),
				.b3(W2L10F),
				.b4(W2L11F),
				.b5(W2L12F),
				.b6(W2L20F),
				.b7(W2L21F),
				.b8(W2L22F),
				.c(c2F00L)
);

assign C200L=c2000L+c2100L+c2200L+c2300L+c2400L+c2500L+c2600L+c2700L+c2800L+c2900L+c2A00L+c2B00L+c2C00L+c2D00L+c2E00L+c2F00L;
assign A200L=(C200L>=0)?1:0;

assign P300L=A200L;

ninexnine_unit ninexnine_unit_6004(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2L000),
				.b1(W2L010),
				.b2(W2L020),
				.b3(W2L100),
				.b4(W2L110),
				.b5(W2L120),
				.b6(W2L200),
				.b7(W2L210),
				.b8(W2L220),
				.c(c2001L)
);

ninexnine_unit ninexnine_unit_6005(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2L001),
				.b1(W2L011),
				.b2(W2L021),
				.b3(W2L101),
				.b4(W2L111),
				.b5(W2L121),
				.b6(W2L201),
				.b7(W2L211),
				.b8(W2L221),
				.c(c2101L)
);

ninexnine_unit ninexnine_unit_6006(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2L002),
				.b1(W2L012),
				.b2(W2L022),
				.b3(W2L102),
				.b4(W2L112),
				.b5(W2L122),
				.b6(W2L202),
				.b7(W2L212),
				.b8(W2L222),
				.c(c2201L)
);

ninexnine_unit ninexnine_unit_6007(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2L003),
				.b1(W2L013),
				.b2(W2L023),
				.b3(W2L103),
				.b4(W2L113),
				.b5(W2L123),
				.b6(W2L203),
				.b7(W2L213),
				.b8(W2L223),
				.c(c2301L)
);

ninexnine_unit ninexnine_unit_6008(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2L004),
				.b1(W2L014),
				.b2(W2L024),
				.b3(W2L104),
				.b4(W2L114),
				.b5(W2L124),
				.b6(W2L204),
				.b7(W2L214),
				.b8(W2L224),
				.c(c2401L)
);

ninexnine_unit ninexnine_unit_6009(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2L005),
				.b1(W2L015),
				.b2(W2L025),
				.b3(W2L105),
				.b4(W2L115),
				.b5(W2L125),
				.b6(W2L205),
				.b7(W2L215),
				.b8(W2L225),
				.c(c2501L)
);

ninexnine_unit ninexnine_unit_6010(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2L006),
				.b1(W2L016),
				.b2(W2L026),
				.b3(W2L106),
				.b4(W2L116),
				.b5(W2L126),
				.b6(W2L206),
				.b7(W2L216),
				.b8(W2L226),
				.c(c2601L)
);

ninexnine_unit ninexnine_unit_6011(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2L007),
				.b1(W2L017),
				.b2(W2L027),
				.b3(W2L107),
				.b4(W2L117),
				.b5(W2L127),
				.b6(W2L207),
				.b7(W2L217),
				.b8(W2L227),
				.c(c2701L)
);

ninexnine_unit ninexnine_unit_6012(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2L008),
				.b1(W2L018),
				.b2(W2L028),
				.b3(W2L108),
				.b4(W2L118),
				.b5(W2L128),
				.b6(W2L208),
				.b7(W2L218),
				.b8(W2L228),
				.c(c2801L)
);

ninexnine_unit ninexnine_unit_6013(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2L009),
				.b1(W2L019),
				.b2(W2L029),
				.b3(W2L109),
				.b4(W2L119),
				.b5(W2L129),
				.b6(W2L209),
				.b7(W2L219),
				.b8(W2L229),
				.c(c2901L)
);

ninexnine_unit ninexnine_unit_6014(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2L00A),
				.b1(W2L01A),
				.b2(W2L02A),
				.b3(W2L10A),
				.b4(W2L11A),
				.b5(W2L12A),
				.b6(W2L20A),
				.b7(W2L21A),
				.b8(W2L22A),
				.c(c2A01L)
);

ninexnine_unit ninexnine_unit_6015(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2L00B),
				.b1(W2L01B),
				.b2(W2L02B),
				.b3(W2L10B),
				.b4(W2L11B),
				.b5(W2L12B),
				.b6(W2L20B),
				.b7(W2L21B),
				.b8(W2L22B),
				.c(c2B01L)
);

ninexnine_unit ninexnine_unit_6016(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2L00C),
				.b1(W2L01C),
				.b2(W2L02C),
				.b3(W2L10C),
				.b4(W2L11C),
				.b5(W2L12C),
				.b6(W2L20C),
				.b7(W2L21C),
				.b8(W2L22C),
				.c(c2C01L)
);

ninexnine_unit ninexnine_unit_6017(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2L00D),
				.b1(W2L01D),
				.b2(W2L02D),
				.b3(W2L10D),
				.b4(W2L11D),
				.b5(W2L12D),
				.b6(W2L20D),
				.b7(W2L21D),
				.b8(W2L22D),
				.c(c2D01L)
);

ninexnine_unit ninexnine_unit_6018(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2L00E),
				.b1(W2L01E),
				.b2(W2L02E),
				.b3(W2L10E),
				.b4(W2L11E),
				.b5(W2L12E),
				.b6(W2L20E),
				.b7(W2L21E),
				.b8(W2L22E),
				.c(c2E01L)
);

ninexnine_unit ninexnine_unit_6019(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2L00F),
				.b1(W2L01F),
				.b2(W2L02F),
				.b3(W2L10F),
				.b4(W2L11F),
				.b5(W2L12F),
				.b6(W2L20F),
				.b7(W2L21F),
				.b8(W2L22F),
				.c(c2F01L)
);

assign C201L=c2001L+c2101L+c2201L+c2301L+c2401L+c2501L+c2601L+c2701L+c2801L+c2901L+c2A01L+c2B01L+c2C01L+c2D01L+c2E01L+c2F01L;
assign A201L=(C201L>=0)?1:0;

assign P301L=A201L;

ninexnine_unit ninexnine_unit_6020(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2L000),
				.b1(W2L010),
				.b2(W2L020),
				.b3(W2L100),
				.b4(W2L110),
				.b5(W2L120),
				.b6(W2L200),
				.b7(W2L210),
				.b8(W2L220),
				.c(c2002L)
);

ninexnine_unit ninexnine_unit_6021(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2L001),
				.b1(W2L011),
				.b2(W2L021),
				.b3(W2L101),
				.b4(W2L111),
				.b5(W2L121),
				.b6(W2L201),
				.b7(W2L211),
				.b8(W2L221),
				.c(c2102L)
);

ninexnine_unit ninexnine_unit_6022(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2L002),
				.b1(W2L012),
				.b2(W2L022),
				.b3(W2L102),
				.b4(W2L112),
				.b5(W2L122),
				.b6(W2L202),
				.b7(W2L212),
				.b8(W2L222),
				.c(c2202L)
);

ninexnine_unit ninexnine_unit_6023(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2L003),
				.b1(W2L013),
				.b2(W2L023),
				.b3(W2L103),
				.b4(W2L113),
				.b5(W2L123),
				.b6(W2L203),
				.b7(W2L213),
				.b8(W2L223),
				.c(c2302L)
);

ninexnine_unit ninexnine_unit_6024(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2L004),
				.b1(W2L014),
				.b2(W2L024),
				.b3(W2L104),
				.b4(W2L114),
				.b5(W2L124),
				.b6(W2L204),
				.b7(W2L214),
				.b8(W2L224),
				.c(c2402L)
);

ninexnine_unit ninexnine_unit_6025(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2L005),
				.b1(W2L015),
				.b2(W2L025),
				.b3(W2L105),
				.b4(W2L115),
				.b5(W2L125),
				.b6(W2L205),
				.b7(W2L215),
				.b8(W2L225),
				.c(c2502L)
);

ninexnine_unit ninexnine_unit_6026(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2L006),
				.b1(W2L016),
				.b2(W2L026),
				.b3(W2L106),
				.b4(W2L116),
				.b5(W2L126),
				.b6(W2L206),
				.b7(W2L216),
				.b8(W2L226),
				.c(c2602L)
);

ninexnine_unit ninexnine_unit_6027(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2L007),
				.b1(W2L017),
				.b2(W2L027),
				.b3(W2L107),
				.b4(W2L117),
				.b5(W2L127),
				.b6(W2L207),
				.b7(W2L217),
				.b8(W2L227),
				.c(c2702L)
);

ninexnine_unit ninexnine_unit_6028(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2L008),
				.b1(W2L018),
				.b2(W2L028),
				.b3(W2L108),
				.b4(W2L118),
				.b5(W2L128),
				.b6(W2L208),
				.b7(W2L218),
				.b8(W2L228),
				.c(c2802L)
);

ninexnine_unit ninexnine_unit_6029(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2L009),
				.b1(W2L019),
				.b2(W2L029),
				.b3(W2L109),
				.b4(W2L119),
				.b5(W2L129),
				.b6(W2L209),
				.b7(W2L219),
				.b8(W2L229),
				.c(c2902L)
);

ninexnine_unit ninexnine_unit_6030(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2L00A),
				.b1(W2L01A),
				.b2(W2L02A),
				.b3(W2L10A),
				.b4(W2L11A),
				.b5(W2L12A),
				.b6(W2L20A),
				.b7(W2L21A),
				.b8(W2L22A),
				.c(c2A02L)
);

ninexnine_unit ninexnine_unit_6031(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2L00B),
				.b1(W2L01B),
				.b2(W2L02B),
				.b3(W2L10B),
				.b4(W2L11B),
				.b5(W2L12B),
				.b6(W2L20B),
				.b7(W2L21B),
				.b8(W2L22B),
				.c(c2B02L)
);

ninexnine_unit ninexnine_unit_6032(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2L00C),
				.b1(W2L01C),
				.b2(W2L02C),
				.b3(W2L10C),
				.b4(W2L11C),
				.b5(W2L12C),
				.b6(W2L20C),
				.b7(W2L21C),
				.b8(W2L22C),
				.c(c2C02L)
);

ninexnine_unit ninexnine_unit_6033(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2L00D),
				.b1(W2L01D),
				.b2(W2L02D),
				.b3(W2L10D),
				.b4(W2L11D),
				.b5(W2L12D),
				.b6(W2L20D),
				.b7(W2L21D),
				.b8(W2L22D),
				.c(c2D02L)
);

ninexnine_unit ninexnine_unit_6034(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2L00E),
				.b1(W2L01E),
				.b2(W2L02E),
				.b3(W2L10E),
				.b4(W2L11E),
				.b5(W2L12E),
				.b6(W2L20E),
				.b7(W2L21E),
				.b8(W2L22E),
				.c(c2E02L)
);

ninexnine_unit ninexnine_unit_6035(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2L00F),
				.b1(W2L01F),
				.b2(W2L02F),
				.b3(W2L10F),
				.b4(W2L11F),
				.b5(W2L12F),
				.b6(W2L20F),
				.b7(W2L21F),
				.b8(W2L22F),
				.c(c2F02L)
);

assign C202L=c2002L+c2102L+c2202L+c2302L+c2402L+c2502L+c2602L+c2702L+c2802L+c2902L+c2A02L+c2B02L+c2C02L+c2D02L+c2E02L+c2F02L;
assign A202L=(C202L>=0)?1:0;

assign P302L=A202L;

ninexnine_unit ninexnine_unit_6036(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2L000),
				.b1(W2L010),
				.b2(W2L020),
				.b3(W2L100),
				.b4(W2L110),
				.b5(W2L120),
				.b6(W2L200),
				.b7(W2L210),
				.b8(W2L220),
				.c(c2010L)
);

ninexnine_unit ninexnine_unit_6037(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2L001),
				.b1(W2L011),
				.b2(W2L021),
				.b3(W2L101),
				.b4(W2L111),
				.b5(W2L121),
				.b6(W2L201),
				.b7(W2L211),
				.b8(W2L221),
				.c(c2110L)
);

ninexnine_unit ninexnine_unit_6038(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2L002),
				.b1(W2L012),
				.b2(W2L022),
				.b3(W2L102),
				.b4(W2L112),
				.b5(W2L122),
				.b6(W2L202),
				.b7(W2L212),
				.b8(W2L222),
				.c(c2210L)
);

ninexnine_unit ninexnine_unit_6039(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2L003),
				.b1(W2L013),
				.b2(W2L023),
				.b3(W2L103),
				.b4(W2L113),
				.b5(W2L123),
				.b6(W2L203),
				.b7(W2L213),
				.b8(W2L223),
				.c(c2310L)
);

ninexnine_unit ninexnine_unit_6040(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2L004),
				.b1(W2L014),
				.b2(W2L024),
				.b3(W2L104),
				.b4(W2L114),
				.b5(W2L124),
				.b6(W2L204),
				.b7(W2L214),
				.b8(W2L224),
				.c(c2410L)
);

ninexnine_unit ninexnine_unit_6041(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2L005),
				.b1(W2L015),
				.b2(W2L025),
				.b3(W2L105),
				.b4(W2L115),
				.b5(W2L125),
				.b6(W2L205),
				.b7(W2L215),
				.b8(W2L225),
				.c(c2510L)
);

ninexnine_unit ninexnine_unit_6042(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2L006),
				.b1(W2L016),
				.b2(W2L026),
				.b3(W2L106),
				.b4(W2L116),
				.b5(W2L126),
				.b6(W2L206),
				.b7(W2L216),
				.b8(W2L226),
				.c(c2610L)
);

ninexnine_unit ninexnine_unit_6043(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2L007),
				.b1(W2L017),
				.b2(W2L027),
				.b3(W2L107),
				.b4(W2L117),
				.b5(W2L127),
				.b6(W2L207),
				.b7(W2L217),
				.b8(W2L227),
				.c(c2710L)
);

ninexnine_unit ninexnine_unit_6044(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2L008),
				.b1(W2L018),
				.b2(W2L028),
				.b3(W2L108),
				.b4(W2L118),
				.b5(W2L128),
				.b6(W2L208),
				.b7(W2L218),
				.b8(W2L228),
				.c(c2810L)
);

ninexnine_unit ninexnine_unit_6045(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2L009),
				.b1(W2L019),
				.b2(W2L029),
				.b3(W2L109),
				.b4(W2L119),
				.b5(W2L129),
				.b6(W2L209),
				.b7(W2L219),
				.b8(W2L229),
				.c(c2910L)
);

ninexnine_unit ninexnine_unit_6046(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2L00A),
				.b1(W2L01A),
				.b2(W2L02A),
				.b3(W2L10A),
				.b4(W2L11A),
				.b5(W2L12A),
				.b6(W2L20A),
				.b7(W2L21A),
				.b8(W2L22A),
				.c(c2A10L)
);

ninexnine_unit ninexnine_unit_6047(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2L00B),
				.b1(W2L01B),
				.b2(W2L02B),
				.b3(W2L10B),
				.b4(W2L11B),
				.b5(W2L12B),
				.b6(W2L20B),
				.b7(W2L21B),
				.b8(W2L22B),
				.c(c2B10L)
);

ninexnine_unit ninexnine_unit_6048(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2L00C),
				.b1(W2L01C),
				.b2(W2L02C),
				.b3(W2L10C),
				.b4(W2L11C),
				.b5(W2L12C),
				.b6(W2L20C),
				.b7(W2L21C),
				.b8(W2L22C),
				.c(c2C10L)
);

ninexnine_unit ninexnine_unit_6049(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2L00D),
				.b1(W2L01D),
				.b2(W2L02D),
				.b3(W2L10D),
				.b4(W2L11D),
				.b5(W2L12D),
				.b6(W2L20D),
				.b7(W2L21D),
				.b8(W2L22D),
				.c(c2D10L)
);

ninexnine_unit ninexnine_unit_6050(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2L00E),
				.b1(W2L01E),
				.b2(W2L02E),
				.b3(W2L10E),
				.b4(W2L11E),
				.b5(W2L12E),
				.b6(W2L20E),
				.b7(W2L21E),
				.b8(W2L22E),
				.c(c2E10L)
);

ninexnine_unit ninexnine_unit_6051(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2L00F),
				.b1(W2L01F),
				.b2(W2L02F),
				.b3(W2L10F),
				.b4(W2L11F),
				.b5(W2L12F),
				.b6(W2L20F),
				.b7(W2L21F),
				.b8(W2L22F),
				.c(c2F10L)
);

assign C210L=c2010L+c2110L+c2210L+c2310L+c2410L+c2510L+c2610L+c2710L+c2810L+c2910L+c2A10L+c2B10L+c2C10L+c2D10L+c2E10L+c2F10L;
assign A210L=(C210L>=0)?1:0;

assign P310L=A210L;

ninexnine_unit ninexnine_unit_6052(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2L000),
				.b1(W2L010),
				.b2(W2L020),
				.b3(W2L100),
				.b4(W2L110),
				.b5(W2L120),
				.b6(W2L200),
				.b7(W2L210),
				.b8(W2L220),
				.c(c2011L)
);

ninexnine_unit ninexnine_unit_6053(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2L001),
				.b1(W2L011),
				.b2(W2L021),
				.b3(W2L101),
				.b4(W2L111),
				.b5(W2L121),
				.b6(W2L201),
				.b7(W2L211),
				.b8(W2L221),
				.c(c2111L)
);

ninexnine_unit ninexnine_unit_6054(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2L002),
				.b1(W2L012),
				.b2(W2L022),
				.b3(W2L102),
				.b4(W2L112),
				.b5(W2L122),
				.b6(W2L202),
				.b7(W2L212),
				.b8(W2L222),
				.c(c2211L)
);

ninexnine_unit ninexnine_unit_6055(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2L003),
				.b1(W2L013),
				.b2(W2L023),
				.b3(W2L103),
				.b4(W2L113),
				.b5(W2L123),
				.b6(W2L203),
				.b7(W2L213),
				.b8(W2L223),
				.c(c2311L)
);

ninexnine_unit ninexnine_unit_6056(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2L004),
				.b1(W2L014),
				.b2(W2L024),
				.b3(W2L104),
				.b4(W2L114),
				.b5(W2L124),
				.b6(W2L204),
				.b7(W2L214),
				.b8(W2L224),
				.c(c2411L)
);

ninexnine_unit ninexnine_unit_6057(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2L005),
				.b1(W2L015),
				.b2(W2L025),
				.b3(W2L105),
				.b4(W2L115),
				.b5(W2L125),
				.b6(W2L205),
				.b7(W2L215),
				.b8(W2L225),
				.c(c2511L)
);

ninexnine_unit ninexnine_unit_6058(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2L006),
				.b1(W2L016),
				.b2(W2L026),
				.b3(W2L106),
				.b4(W2L116),
				.b5(W2L126),
				.b6(W2L206),
				.b7(W2L216),
				.b8(W2L226),
				.c(c2611L)
);

ninexnine_unit ninexnine_unit_6059(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2L007),
				.b1(W2L017),
				.b2(W2L027),
				.b3(W2L107),
				.b4(W2L117),
				.b5(W2L127),
				.b6(W2L207),
				.b7(W2L217),
				.b8(W2L227),
				.c(c2711L)
);

ninexnine_unit ninexnine_unit_6060(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2L008),
				.b1(W2L018),
				.b2(W2L028),
				.b3(W2L108),
				.b4(W2L118),
				.b5(W2L128),
				.b6(W2L208),
				.b7(W2L218),
				.b8(W2L228),
				.c(c2811L)
);

ninexnine_unit ninexnine_unit_6061(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2L009),
				.b1(W2L019),
				.b2(W2L029),
				.b3(W2L109),
				.b4(W2L119),
				.b5(W2L129),
				.b6(W2L209),
				.b7(W2L219),
				.b8(W2L229),
				.c(c2911L)
);

ninexnine_unit ninexnine_unit_6062(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2L00A),
				.b1(W2L01A),
				.b2(W2L02A),
				.b3(W2L10A),
				.b4(W2L11A),
				.b5(W2L12A),
				.b6(W2L20A),
				.b7(W2L21A),
				.b8(W2L22A),
				.c(c2A11L)
);

ninexnine_unit ninexnine_unit_6063(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2L00B),
				.b1(W2L01B),
				.b2(W2L02B),
				.b3(W2L10B),
				.b4(W2L11B),
				.b5(W2L12B),
				.b6(W2L20B),
				.b7(W2L21B),
				.b8(W2L22B),
				.c(c2B11L)
);

ninexnine_unit ninexnine_unit_6064(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2L00C),
				.b1(W2L01C),
				.b2(W2L02C),
				.b3(W2L10C),
				.b4(W2L11C),
				.b5(W2L12C),
				.b6(W2L20C),
				.b7(W2L21C),
				.b8(W2L22C),
				.c(c2C11L)
);

ninexnine_unit ninexnine_unit_6065(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2L00D),
				.b1(W2L01D),
				.b2(W2L02D),
				.b3(W2L10D),
				.b4(W2L11D),
				.b5(W2L12D),
				.b6(W2L20D),
				.b7(W2L21D),
				.b8(W2L22D),
				.c(c2D11L)
);

ninexnine_unit ninexnine_unit_6066(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2L00E),
				.b1(W2L01E),
				.b2(W2L02E),
				.b3(W2L10E),
				.b4(W2L11E),
				.b5(W2L12E),
				.b6(W2L20E),
				.b7(W2L21E),
				.b8(W2L22E),
				.c(c2E11L)
);

ninexnine_unit ninexnine_unit_6067(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2L00F),
				.b1(W2L01F),
				.b2(W2L02F),
				.b3(W2L10F),
				.b4(W2L11F),
				.b5(W2L12F),
				.b6(W2L20F),
				.b7(W2L21F),
				.b8(W2L22F),
				.c(c2F11L)
);

assign C211L=c2011L+c2111L+c2211L+c2311L+c2411L+c2511L+c2611L+c2711L+c2811L+c2911L+c2A11L+c2B11L+c2C11L+c2D11L+c2E11L+c2F11L;
assign A211L=(C211L>=0)?1:0;

assign P311L=A211L;

ninexnine_unit ninexnine_unit_6068(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2L000),
				.b1(W2L010),
				.b2(W2L020),
				.b3(W2L100),
				.b4(W2L110),
				.b5(W2L120),
				.b6(W2L200),
				.b7(W2L210),
				.b8(W2L220),
				.c(c2012L)
);

ninexnine_unit ninexnine_unit_6069(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2L001),
				.b1(W2L011),
				.b2(W2L021),
				.b3(W2L101),
				.b4(W2L111),
				.b5(W2L121),
				.b6(W2L201),
				.b7(W2L211),
				.b8(W2L221),
				.c(c2112L)
);

ninexnine_unit ninexnine_unit_6070(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2L002),
				.b1(W2L012),
				.b2(W2L022),
				.b3(W2L102),
				.b4(W2L112),
				.b5(W2L122),
				.b6(W2L202),
				.b7(W2L212),
				.b8(W2L222),
				.c(c2212L)
);

ninexnine_unit ninexnine_unit_6071(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2L003),
				.b1(W2L013),
				.b2(W2L023),
				.b3(W2L103),
				.b4(W2L113),
				.b5(W2L123),
				.b6(W2L203),
				.b7(W2L213),
				.b8(W2L223),
				.c(c2312L)
);

ninexnine_unit ninexnine_unit_6072(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2L004),
				.b1(W2L014),
				.b2(W2L024),
				.b3(W2L104),
				.b4(W2L114),
				.b5(W2L124),
				.b6(W2L204),
				.b7(W2L214),
				.b8(W2L224),
				.c(c2412L)
);

ninexnine_unit ninexnine_unit_6073(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2L005),
				.b1(W2L015),
				.b2(W2L025),
				.b3(W2L105),
				.b4(W2L115),
				.b5(W2L125),
				.b6(W2L205),
				.b7(W2L215),
				.b8(W2L225),
				.c(c2512L)
);

ninexnine_unit ninexnine_unit_6074(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2L006),
				.b1(W2L016),
				.b2(W2L026),
				.b3(W2L106),
				.b4(W2L116),
				.b5(W2L126),
				.b6(W2L206),
				.b7(W2L216),
				.b8(W2L226),
				.c(c2612L)
);

ninexnine_unit ninexnine_unit_6075(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2L007),
				.b1(W2L017),
				.b2(W2L027),
				.b3(W2L107),
				.b4(W2L117),
				.b5(W2L127),
				.b6(W2L207),
				.b7(W2L217),
				.b8(W2L227),
				.c(c2712L)
);

ninexnine_unit ninexnine_unit_6076(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2L008),
				.b1(W2L018),
				.b2(W2L028),
				.b3(W2L108),
				.b4(W2L118),
				.b5(W2L128),
				.b6(W2L208),
				.b7(W2L218),
				.b8(W2L228),
				.c(c2812L)
);

ninexnine_unit ninexnine_unit_6077(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2L009),
				.b1(W2L019),
				.b2(W2L029),
				.b3(W2L109),
				.b4(W2L119),
				.b5(W2L129),
				.b6(W2L209),
				.b7(W2L219),
				.b8(W2L229),
				.c(c2912L)
);

ninexnine_unit ninexnine_unit_6078(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2L00A),
				.b1(W2L01A),
				.b2(W2L02A),
				.b3(W2L10A),
				.b4(W2L11A),
				.b5(W2L12A),
				.b6(W2L20A),
				.b7(W2L21A),
				.b8(W2L22A),
				.c(c2A12L)
);

ninexnine_unit ninexnine_unit_6079(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2L00B),
				.b1(W2L01B),
				.b2(W2L02B),
				.b3(W2L10B),
				.b4(W2L11B),
				.b5(W2L12B),
				.b6(W2L20B),
				.b7(W2L21B),
				.b8(W2L22B),
				.c(c2B12L)
);

ninexnine_unit ninexnine_unit_6080(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2L00C),
				.b1(W2L01C),
				.b2(W2L02C),
				.b3(W2L10C),
				.b4(W2L11C),
				.b5(W2L12C),
				.b6(W2L20C),
				.b7(W2L21C),
				.b8(W2L22C),
				.c(c2C12L)
);

ninexnine_unit ninexnine_unit_6081(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2L00D),
				.b1(W2L01D),
				.b2(W2L02D),
				.b3(W2L10D),
				.b4(W2L11D),
				.b5(W2L12D),
				.b6(W2L20D),
				.b7(W2L21D),
				.b8(W2L22D),
				.c(c2D12L)
);

ninexnine_unit ninexnine_unit_6082(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2L00E),
				.b1(W2L01E),
				.b2(W2L02E),
				.b3(W2L10E),
				.b4(W2L11E),
				.b5(W2L12E),
				.b6(W2L20E),
				.b7(W2L21E),
				.b8(W2L22E),
				.c(c2E12L)
);

ninexnine_unit ninexnine_unit_6083(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2L00F),
				.b1(W2L01F),
				.b2(W2L02F),
				.b3(W2L10F),
				.b4(W2L11F),
				.b5(W2L12F),
				.b6(W2L20F),
				.b7(W2L21F),
				.b8(W2L22F),
				.c(c2F12L)
);

assign C212L=c2012L+c2112L+c2212L+c2312L+c2412L+c2512L+c2612L+c2712L+c2812L+c2912L+c2A12L+c2B12L+c2C12L+c2D12L+c2E12L+c2F12L;
assign A212L=(C212L>=0)?1:0;

assign P312L=A212L;

ninexnine_unit ninexnine_unit_6084(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2L000),
				.b1(W2L010),
				.b2(W2L020),
				.b3(W2L100),
				.b4(W2L110),
				.b5(W2L120),
				.b6(W2L200),
				.b7(W2L210),
				.b8(W2L220),
				.c(c2020L)
);

ninexnine_unit ninexnine_unit_6085(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2L001),
				.b1(W2L011),
				.b2(W2L021),
				.b3(W2L101),
				.b4(W2L111),
				.b5(W2L121),
				.b6(W2L201),
				.b7(W2L211),
				.b8(W2L221),
				.c(c2120L)
);

ninexnine_unit ninexnine_unit_6086(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2L002),
				.b1(W2L012),
				.b2(W2L022),
				.b3(W2L102),
				.b4(W2L112),
				.b5(W2L122),
				.b6(W2L202),
				.b7(W2L212),
				.b8(W2L222),
				.c(c2220L)
);

ninexnine_unit ninexnine_unit_6087(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2L003),
				.b1(W2L013),
				.b2(W2L023),
				.b3(W2L103),
				.b4(W2L113),
				.b5(W2L123),
				.b6(W2L203),
				.b7(W2L213),
				.b8(W2L223),
				.c(c2320L)
);

ninexnine_unit ninexnine_unit_6088(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2L004),
				.b1(W2L014),
				.b2(W2L024),
				.b3(W2L104),
				.b4(W2L114),
				.b5(W2L124),
				.b6(W2L204),
				.b7(W2L214),
				.b8(W2L224),
				.c(c2420L)
);

ninexnine_unit ninexnine_unit_6089(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2L005),
				.b1(W2L015),
				.b2(W2L025),
				.b3(W2L105),
				.b4(W2L115),
				.b5(W2L125),
				.b6(W2L205),
				.b7(W2L215),
				.b8(W2L225),
				.c(c2520L)
);

ninexnine_unit ninexnine_unit_6090(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2L006),
				.b1(W2L016),
				.b2(W2L026),
				.b3(W2L106),
				.b4(W2L116),
				.b5(W2L126),
				.b6(W2L206),
				.b7(W2L216),
				.b8(W2L226),
				.c(c2620L)
);

ninexnine_unit ninexnine_unit_6091(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2L007),
				.b1(W2L017),
				.b2(W2L027),
				.b3(W2L107),
				.b4(W2L117),
				.b5(W2L127),
				.b6(W2L207),
				.b7(W2L217),
				.b8(W2L227),
				.c(c2720L)
);

ninexnine_unit ninexnine_unit_6092(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2L008),
				.b1(W2L018),
				.b2(W2L028),
				.b3(W2L108),
				.b4(W2L118),
				.b5(W2L128),
				.b6(W2L208),
				.b7(W2L218),
				.b8(W2L228),
				.c(c2820L)
);

ninexnine_unit ninexnine_unit_6093(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2L009),
				.b1(W2L019),
				.b2(W2L029),
				.b3(W2L109),
				.b4(W2L119),
				.b5(W2L129),
				.b6(W2L209),
				.b7(W2L219),
				.b8(W2L229),
				.c(c2920L)
);

ninexnine_unit ninexnine_unit_6094(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2L00A),
				.b1(W2L01A),
				.b2(W2L02A),
				.b3(W2L10A),
				.b4(W2L11A),
				.b5(W2L12A),
				.b6(W2L20A),
				.b7(W2L21A),
				.b8(W2L22A),
				.c(c2A20L)
);

ninexnine_unit ninexnine_unit_6095(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2L00B),
				.b1(W2L01B),
				.b2(W2L02B),
				.b3(W2L10B),
				.b4(W2L11B),
				.b5(W2L12B),
				.b6(W2L20B),
				.b7(W2L21B),
				.b8(W2L22B),
				.c(c2B20L)
);

ninexnine_unit ninexnine_unit_6096(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2L00C),
				.b1(W2L01C),
				.b2(W2L02C),
				.b3(W2L10C),
				.b4(W2L11C),
				.b5(W2L12C),
				.b6(W2L20C),
				.b7(W2L21C),
				.b8(W2L22C),
				.c(c2C20L)
);

ninexnine_unit ninexnine_unit_6097(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2L00D),
				.b1(W2L01D),
				.b2(W2L02D),
				.b3(W2L10D),
				.b4(W2L11D),
				.b5(W2L12D),
				.b6(W2L20D),
				.b7(W2L21D),
				.b8(W2L22D),
				.c(c2D20L)
);

ninexnine_unit ninexnine_unit_6098(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2L00E),
				.b1(W2L01E),
				.b2(W2L02E),
				.b3(W2L10E),
				.b4(W2L11E),
				.b5(W2L12E),
				.b6(W2L20E),
				.b7(W2L21E),
				.b8(W2L22E),
				.c(c2E20L)
);

ninexnine_unit ninexnine_unit_6099(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2L00F),
				.b1(W2L01F),
				.b2(W2L02F),
				.b3(W2L10F),
				.b4(W2L11F),
				.b5(W2L12F),
				.b6(W2L20F),
				.b7(W2L21F),
				.b8(W2L22F),
				.c(c2F20L)
);

assign C220L=c2020L+c2120L+c2220L+c2320L+c2420L+c2520L+c2620L+c2720L+c2820L+c2920L+c2A20L+c2B20L+c2C20L+c2D20L+c2E20L+c2F20L;
assign A220L=(C220L>=0)?1:0;

assign P320L=A220L;

ninexnine_unit ninexnine_unit_6100(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2L000),
				.b1(W2L010),
				.b2(W2L020),
				.b3(W2L100),
				.b4(W2L110),
				.b5(W2L120),
				.b6(W2L200),
				.b7(W2L210),
				.b8(W2L220),
				.c(c2021L)
);

ninexnine_unit ninexnine_unit_6101(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2L001),
				.b1(W2L011),
				.b2(W2L021),
				.b3(W2L101),
				.b4(W2L111),
				.b5(W2L121),
				.b6(W2L201),
				.b7(W2L211),
				.b8(W2L221),
				.c(c2121L)
);

ninexnine_unit ninexnine_unit_6102(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2L002),
				.b1(W2L012),
				.b2(W2L022),
				.b3(W2L102),
				.b4(W2L112),
				.b5(W2L122),
				.b6(W2L202),
				.b7(W2L212),
				.b8(W2L222),
				.c(c2221L)
);

ninexnine_unit ninexnine_unit_6103(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2L003),
				.b1(W2L013),
				.b2(W2L023),
				.b3(W2L103),
				.b4(W2L113),
				.b5(W2L123),
				.b6(W2L203),
				.b7(W2L213),
				.b8(W2L223),
				.c(c2321L)
);

ninexnine_unit ninexnine_unit_6104(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2L004),
				.b1(W2L014),
				.b2(W2L024),
				.b3(W2L104),
				.b4(W2L114),
				.b5(W2L124),
				.b6(W2L204),
				.b7(W2L214),
				.b8(W2L224),
				.c(c2421L)
);

ninexnine_unit ninexnine_unit_6105(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2L005),
				.b1(W2L015),
				.b2(W2L025),
				.b3(W2L105),
				.b4(W2L115),
				.b5(W2L125),
				.b6(W2L205),
				.b7(W2L215),
				.b8(W2L225),
				.c(c2521L)
);

ninexnine_unit ninexnine_unit_6106(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2L006),
				.b1(W2L016),
				.b2(W2L026),
				.b3(W2L106),
				.b4(W2L116),
				.b5(W2L126),
				.b6(W2L206),
				.b7(W2L216),
				.b8(W2L226),
				.c(c2621L)
);

ninexnine_unit ninexnine_unit_6107(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2L007),
				.b1(W2L017),
				.b2(W2L027),
				.b3(W2L107),
				.b4(W2L117),
				.b5(W2L127),
				.b6(W2L207),
				.b7(W2L217),
				.b8(W2L227),
				.c(c2721L)
);

ninexnine_unit ninexnine_unit_6108(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2L008),
				.b1(W2L018),
				.b2(W2L028),
				.b3(W2L108),
				.b4(W2L118),
				.b5(W2L128),
				.b6(W2L208),
				.b7(W2L218),
				.b8(W2L228),
				.c(c2821L)
);

ninexnine_unit ninexnine_unit_6109(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2L009),
				.b1(W2L019),
				.b2(W2L029),
				.b3(W2L109),
				.b4(W2L119),
				.b5(W2L129),
				.b6(W2L209),
				.b7(W2L219),
				.b8(W2L229),
				.c(c2921L)
);

ninexnine_unit ninexnine_unit_6110(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2L00A),
				.b1(W2L01A),
				.b2(W2L02A),
				.b3(W2L10A),
				.b4(W2L11A),
				.b5(W2L12A),
				.b6(W2L20A),
				.b7(W2L21A),
				.b8(W2L22A),
				.c(c2A21L)
);

ninexnine_unit ninexnine_unit_6111(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2L00B),
				.b1(W2L01B),
				.b2(W2L02B),
				.b3(W2L10B),
				.b4(W2L11B),
				.b5(W2L12B),
				.b6(W2L20B),
				.b7(W2L21B),
				.b8(W2L22B),
				.c(c2B21L)
);

ninexnine_unit ninexnine_unit_6112(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2L00C),
				.b1(W2L01C),
				.b2(W2L02C),
				.b3(W2L10C),
				.b4(W2L11C),
				.b5(W2L12C),
				.b6(W2L20C),
				.b7(W2L21C),
				.b8(W2L22C),
				.c(c2C21L)
);

ninexnine_unit ninexnine_unit_6113(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2L00D),
				.b1(W2L01D),
				.b2(W2L02D),
				.b3(W2L10D),
				.b4(W2L11D),
				.b5(W2L12D),
				.b6(W2L20D),
				.b7(W2L21D),
				.b8(W2L22D),
				.c(c2D21L)
);

ninexnine_unit ninexnine_unit_6114(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2L00E),
				.b1(W2L01E),
				.b2(W2L02E),
				.b3(W2L10E),
				.b4(W2L11E),
				.b5(W2L12E),
				.b6(W2L20E),
				.b7(W2L21E),
				.b8(W2L22E),
				.c(c2E21L)
);

ninexnine_unit ninexnine_unit_6115(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2L00F),
				.b1(W2L01F),
				.b2(W2L02F),
				.b3(W2L10F),
				.b4(W2L11F),
				.b5(W2L12F),
				.b6(W2L20F),
				.b7(W2L21F),
				.b8(W2L22F),
				.c(c2F21L)
);

assign C221L=c2021L+c2121L+c2221L+c2321L+c2421L+c2521L+c2621L+c2721L+c2821L+c2921L+c2A21L+c2B21L+c2C21L+c2D21L+c2E21L+c2F21L;
assign A221L=(C221L>=0)?1:0;

assign P321L=A221L;

ninexnine_unit ninexnine_unit_6116(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2L000),
				.b1(W2L010),
				.b2(W2L020),
				.b3(W2L100),
				.b4(W2L110),
				.b5(W2L120),
				.b6(W2L200),
				.b7(W2L210),
				.b8(W2L220),
				.c(c2022L)
);

ninexnine_unit ninexnine_unit_6117(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2L001),
				.b1(W2L011),
				.b2(W2L021),
				.b3(W2L101),
				.b4(W2L111),
				.b5(W2L121),
				.b6(W2L201),
				.b7(W2L211),
				.b8(W2L221),
				.c(c2122L)
);

ninexnine_unit ninexnine_unit_6118(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2L002),
				.b1(W2L012),
				.b2(W2L022),
				.b3(W2L102),
				.b4(W2L112),
				.b5(W2L122),
				.b6(W2L202),
				.b7(W2L212),
				.b8(W2L222),
				.c(c2222L)
);

ninexnine_unit ninexnine_unit_6119(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2L003),
				.b1(W2L013),
				.b2(W2L023),
				.b3(W2L103),
				.b4(W2L113),
				.b5(W2L123),
				.b6(W2L203),
				.b7(W2L213),
				.b8(W2L223),
				.c(c2322L)
);

ninexnine_unit ninexnine_unit_6120(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2L004),
				.b1(W2L014),
				.b2(W2L024),
				.b3(W2L104),
				.b4(W2L114),
				.b5(W2L124),
				.b6(W2L204),
				.b7(W2L214),
				.b8(W2L224),
				.c(c2422L)
);

ninexnine_unit ninexnine_unit_6121(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2L005),
				.b1(W2L015),
				.b2(W2L025),
				.b3(W2L105),
				.b4(W2L115),
				.b5(W2L125),
				.b6(W2L205),
				.b7(W2L215),
				.b8(W2L225),
				.c(c2522L)
);

ninexnine_unit ninexnine_unit_6122(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2L006),
				.b1(W2L016),
				.b2(W2L026),
				.b3(W2L106),
				.b4(W2L116),
				.b5(W2L126),
				.b6(W2L206),
				.b7(W2L216),
				.b8(W2L226),
				.c(c2622L)
);

ninexnine_unit ninexnine_unit_6123(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2L007),
				.b1(W2L017),
				.b2(W2L027),
				.b3(W2L107),
				.b4(W2L117),
				.b5(W2L127),
				.b6(W2L207),
				.b7(W2L217),
				.b8(W2L227),
				.c(c2722L)
);

ninexnine_unit ninexnine_unit_6124(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2L008),
				.b1(W2L018),
				.b2(W2L028),
				.b3(W2L108),
				.b4(W2L118),
				.b5(W2L128),
				.b6(W2L208),
				.b7(W2L218),
				.b8(W2L228),
				.c(c2822L)
);

ninexnine_unit ninexnine_unit_6125(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2L009),
				.b1(W2L019),
				.b2(W2L029),
				.b3(W2L109),
				.b4(W2L119),
				.b5(W2L129),
				.b6(W2L209),
				.b7(W2L219),
				.b8(W2L229),
				.c(c2922L)
);

ninexnine_unit ninexnine_unit_6126(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2L00A),
				.b1(W2L01A),
				.b2(W2L02A),
				.b3(W2L10A),
				.b4(W2L11A),
				.b5(W2L12A),
				.b6(W2L20A),
				.b7(W2L21A),
				.b8(W2L22A),
				.c(c2A22L)
);

ninexnine_unit ninexnine_unit_6127(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2L00B),
				.b1(W2L01B),
				.b2(W2L02B),
				.b3(W2L10B),
				.b4(W2L11B),
				.b5(W2L12B),
				.b6(W2L20B),
				.b7(W2L21B),
				.b8(W2L22B),
				.c(c2B22L)
);

ninexnine_unit ninexnine_unit_6128(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2L00C),
				.b1(W2L01C),
				.b2(W2L02C),
				.b3(W2L10C),
				.b4(W2L11C),
				.b5(W2L12C),
				.b6(W2L20C),
				.b7(W2L21C),
				.b8(W2L22C),
				.c(c2C22L)
);

ninexnine_unit ninexnine_unit_6129(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2L00D),
				.b1(W2L01D),
				.b2(W2L02D),
				.b3(W2L10D),
				.b4(W2L11D),
				.b5(W2L12D),
				.b6(W2L20D),
				.b7(W2L21D),
				.b8(W2L22D),
				.c(c2D22L)
);

ninexnine_unit ninexnine_unit_6130(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2L00E),
				.b1(W2L01E),
				.b2(W2L02E),
				.b3(W2L10E),
				.b4(W2L11E),
				.b5(W2L12E),
				.b6(W2L20E),
				.b7(W2L21E),
				.b8(W2L22E),
				.c(c2E22L)
);

ninexnine_unit ninexnine_unit_6131(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2L00F),
				.b1(W2L01F),
				.b2(W2L02F),
				.b3(W2L10F),
				.b4(W2L11F),
				.b5(W2L12F),
				.b6(W2L20F),
				.b7(W2L21F),
				.b8(W2L22F),
				.c(c2F22L)
);

assign C222L=c2022L+c2122L+c2222L+c2322L+c2422L+c2522L+c2622L+c2722L+c2822L+c2922L+c2A22L+c2B22L+c2C22L+c2D22L+c2E22L+c2F22L;
assign A222L=(C222L>=0)?1:0;

assign P322L=A222L;

ninexnine_unit ninexnine_unit_6132(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2M000),
				.b1(W2M010),
				.b2(W2M020),
				.b3(W2M100),
				.b4(W2M110),
				.b5(W2M120),
				.b6(W2M200),
				.b7(W2M210),
				.b8(W2M220),
				.c(c2000M)
);

ninexnine_unit ninexnine_unit_6133(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2M001),
				.b1(W2M011),
				.b2(W2M021),
				.b3(W2M101),
				.b4(W2M111),
				.b5(W2M121),
				.b6(W2M201),
				.b7(W2M211),
				.b8(W2M221),
				.c(c2100M)
);

ninexnine_unit ninexnine_unit_6134(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2M002),
				.b1(W2M012),
				.b2(W2M022),
				.b3(W2M102),
				.b4(W2M112),
				.b5(W2M122),
				.b6(W2M202),
				.b7(W2M212),
				.b8(W2M222),
				.c(c2200M)
);

ninexnine_unit ninexnine_unit_6135(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2M003),
				.b1(W2M013),
				.b2(W2M023),
				.b3(W2M103),
				.b4(W2M113),
				.b5(W2M123),
				.b6(W2M203),
				.b7(W2M213),
				.b8(W2M223),
				.c(c2300M)
);

ninexnine_unit ninexnine_unit_6136(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2M004),
				.b1(W2M014),
				.b2(W2M024),
				.b3(W2M104),
				.b4(W2M114),
				.b5(W2M124),
				.b6(W2M204),
				.b7(W2M214),
				.b8(W2M224),
				.c(c2400M)
);

ninexnine_unit ninexnine_unit_6137(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2M005),
				.b1(W2M015),
				.b2(W2M025),
				.b3(W2M105),
				.b4(W2M115),
				.b5(W2M125),
				.b6(W2M205),
				.b7(W2M215),
				.b8(W2M225),
				.c(c2500M)
);

ninexnine_unit ninexnine_unit_6138(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2M006),
				.b1(W2M016),
				.b2(W2M026),
				.b3(W2M106),
				.b4(W2M116),
				.b5(W2M126),
				.b6(W2M206),
				.b7(W2M216),
				.b8(W2M226),
				.c(c2600M)
);

ninexnine_unit ninexnine_unit_6139(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2M007),
				.b1(W2M017),
				.b2(W2M027),
				.b3(W2M107),
				.b4(W2M117),
				.b5(W2M127),
				.b6(W2M207),
				.b7(W2M217),
				.b8(W2M227),
				.c(c2700M)
);

ninexnine_unit ninexnine_unit_6140(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2M008),
				.b1(W2M018),
				.b2(W2M028),
				.b3(W2M108),
				.b4(W2M118),
				.b5(W2M128),
				.b6(W2M208),
				.b7(W2M218),
				.b8(W2M228),
				.c(c2800M)
);

ninexnine_unit ninexnine_unit_6141(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2M009),
				.b1(W2M019),
				.b2(W2M029),
				.b3(W2M109),
				.b4(W2M119),
				.b5(W2M129),
				.b6(W2M209),
				.b7(W2M219),
				.b8(W2M229),
				.c(c2900M)
);

ninexnine_unit ninexnine_unit_6142(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2M00A),
				.b1(W2M01A),
				.b2(W2M02A),
				.b3(W2M10A),
				.b4(W2M11A),
				.b5(W2M12A),
				.b6(W2M20A),
				.b7(W2M21A),
				.b8(W2M22A),
				.c(c2A00M)
);

ninexnine_unit ninexnine_unit_6143(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2M00B),
				.b1(W2M01B),
				.b2(W2M02B),
				.b3(W2M10B),
				.b4(W2M11B),
				.b5(W2M12B),
				.b6(W2M20B),
				.b7(W2M21B),
				.b8(W2M22B),
				.c(c2B00M)
);

ninexnine_unit ninexnine_unit_6144(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2M00C),
				.b1(W2M01C),
				.b2(W2M02C),
				.b3(W2M10C),
				.b4(W2M11C),
				.b5(W2M12C),
				.b6(W2M20C),
				.b7(W2M21C),
				.b8(W2M22C),
				.c(c2C00M)
);

ninexnine_unit ninexnine_unit_6145(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2M00D),
				.b1(W2M01D),
				.b2(W2M02D),
				.b3(W2M10D),
				.b4(W2M11D),
				.b5(W2M12D),
				.b6(W2M20D),
				.b7(W2M21D),
				.b8(W2M22D),
				.c(c2D00M)
);

ninexnine_unit ninexnine_unit_6146(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2M00E),
				.b1(W2M01E),
				.b2(W2M02E),
				.b3(W2M10E),
				.b4(W2M11E),
				.b5(W2M12E),
				.b6(W2M20E),
				.b7(W2M21E),
				.b8(W2M22E),
				.c(c2E00M)
);

ninexnine_unit ninexnine_unit_6147(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2M00F),
				.b1(W2M01F),
				.b2(W2M02F),
				.b3(W2M10F),
				.b4(W2M11F),
				.b5(W2M12F),
				.b6(W2M20F),
				.b7(W2M21F),
				.b8(W2M22F),
				.c(c2F00M)
);

assign C200M=c2000M+c2100M+c2200M+c2300M+c2400M+c2500M+c2600M+c2700M+c2800M+c2900M+c2A00M+c2B00M+c2C00M+c2D00M+c2E00M+c2F00M;
assign A200M=(C200M>=0)?1:0;

assign P300M=A200M;

ninexnine_unit ninexnine_unit_6148(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2M000),
				.b1(W2M010),
				.b2(W2M020),
				.b3(W2M100),
				.b4(W2M110),
				.b5(W2M120),
				.b6(W2M200),
				.b7(W2M210),
				.b8(W2M220),
				.c(c2001M)
);

ninexnine_unit ninexnine_unit_6149(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2M001),
				.b1(W2M011),
				.b2(W2M021),
				.b3(W2M101),
				.b4(W2M111),
				.b5(W2M121),
				.b6(W2M201),
				.b7(W2M211),
				.b8(W2M221),
				.c(c2101M)
);

ninexnine_unit ninexnine_unit_6150(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2M002),
				.b1(W2M012),
				.b2(W2M022),
				.b3(W2M102),
				.b4(W2M112),
				.b5(W2M122),
				.b6(W2M202),
				.b7(W2M212),
				.b8(W2M222),
				.c(c2201M)
);

ninexnine_unit ninexnine_unit_6151(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2M003),
				.b1(W2M013),
				.b2(W2M023),
				.b3(W2M103),
				.b4(W2M113),
				.b5(W2M123),
				.b6(W2M203),
				.b7(W2M213),
				.b8(W2M223),
				.c(c2301M)
);

ninexnine_unit ninexnine_unit_6152(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2M004),
				.b1(W2M014),
				.b2(W2M024),
				.b3(W2M104),
				.b4(W2M114),
				.b5(W2M124),
				.b6(W2M204),
				.b7(W2M214),
				.b8(W2M224),
				.c(c2401M)
);

ninexnine_unit ninexnine_unit_6153(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2M005),
				.b1(W2M015),
				.b2(W2M025),
				.b3(W2M105),
				.b4(W2M115),
				.b5(W2M125),
				.b6(W2M205),
				.b7(W2M215),
				.b8(W2M225),
				.c(c2501M)
);

ninexnine_unit ninexnine_unit_6154(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2M006),
				.b1(W2M016),
				.b2(W2M026),
				.b3(W2M106),
				.b4(W2M116),
				.b5(W2M126),
				.b6(W2M206),
				.b7(W2M216),
				.b8(W2M226),
				.c(c2601M)
);

ninexnine_unit ninexnine_unit_6155(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2M007),
				.b1(W2M017),
				.b2(W2M027),
				.b3(W2M107),
				.b4(W2M117),
				.b5(W2M127),
				.b6(W2M207),
				.b7(W2M217),
				.b8(W2M227),
				.c(c2701M)
);

ninexnine_unit ninexnine_unit_6156(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2M008),
				.b1(W2M018),
				.b2(W2M028),
				.b3(W2M108),
				.b4(W2M118),
				.b5(W2M128),
				.b6(W2M208),
				.b7(W2M218),
				.b8(W2M228),
				.c(c2801M)
);

ninexnine_unit ninexnine_unit_6157(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2M009),
				.b1(W2M019),
				.b2(W2M029),
				.b3(W2M109),
				.b4(W2M119),
				.b5(W2M129),
				.b6(W2M209),
				.b7(W2M219),
				.b8(W2M229),
				.c(c2901M)
);

ninexnine_unit ninexnine_unit_6158(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2M00A),
				.b1(W2M01A),
				.b2(W2M02A),
				.b3(W2M10A),
				.b4(W2M11A),
				.b5(W2M12A),
				.b6(W2M20A),
				.b7(W2M21A),
				.b8(W2M22A),
				.c(c2A01M)
);

ninexnine_unit ninexnine_unit_6159(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2M00B),
				.b1(W2M01B),
				.b2(W2M02B),
				.b3(W2M10B),
				.b4(W2M11B),
				.b5(W2M12B),
				.b6(W2M20B),
				.b7(W2M21B),
				.b8(W2M22B),
				.c(c2B01M)
);

ninexnine_unit ninexnine_unit_6160(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2M00C),
				.b1(W2M01C),
				.b2(W2M02C),
				.b3(W2M10C),
				.b4(W2M11C),
				.b5(W2M12C),
				.b6(W2M20C),
				.b7(W2M21C),
				.b8(W2M22C),
				.c(c2C01M)
);

ninexnine_unit ninexnine_unit_6161(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2M00D),
				.b1(W2M01D),
				.b2(W2M02D),
				.b3(W2M10D),
				.b4(W2M11D),
				.b5(W2M12D),
				.b6(W2M20D),
				.b7(W2M21D),
				.b8(W2M22D),
				.c(c2D01M)
);

ninexnine_unit ninexnine_unit_6162(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2M00E),
				.b1(W2M01E),
				.b2(W2M02E),
				.b3(W2M10E),
				.b4(W2M11E),
				.b5(W2M12E),
				.b6(W2M20E),
				.b7(W2M21E),
				.b8(W2M22E),
				.c(c2E01M)
);

ninexnine_unit ninexnine_unit_6163(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2M00F),
				.b1(W2M01F),
				.b2(W2M02F),
				.b3(W2M10F),
				.b4(W2M11F),
				.b5(W2M12F),
				.b6(W2M20F),
				.b7(W2M21F),
				.b8(W2M22F),
				.c(c2F01M)
);

assign C201M=c2001M+c2101M+c2201M+c2301M+c2401M+c2501M+c2601M+c2701M+c2801M+c2901M+c2A01M+c2B01M+c2C01M+c2D01M+c2E01M+c2F01M;
assign A201M=(C201M>=0)?1:0;

assign P301M=A201M;

ninexnine_unit ninexnine_unit_6164(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2M000),
				.b1(W2M010),
				.b2(W2M020),
				.b3(W2M100),
				.b4(W2M110),
				.b5(W2M120),
				.b6(W2M200),
				.b7(W2M210),
				.b8(W2M220),
				.c(c2002M)
);

ninexnine_unit ninexnine_unit_6165(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2M001),
				.b1(W2M011),
				.b2(W2M021),
				.b3(W2M101),
				.b4(W2M111),
				.b5(W2M121),
				.b6(W2M201),
				.b7(W2M211),
				.b8(W2M221),
				.c(c2102M)
);

ninexnine_unit ninexnine_unit_6166(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2M002),
				.b1(W2M012),
				.b2(W2M022),
				.b3(W2M102),
				.b4(W2M112),
				.b5(W2M122),
				.b6(W2M202),
				.b7(W2M212),
				.b8(W2M222),
				.c(c2202M)
);

ninexnine_unit ninexnine_unit_6167(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2M003),
				.b1(W2M013),
				.b2(W2M023),
				.b3(W2M103),
				.b4(W2M113),
				.b5(W2M123),
				.b6(W2M203),
				.b7(W2M213),
				.b8(W2M223),
				.c(c2302M)
);

ninexnine_unit ninexnine_unit_6168(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2M004),
				.b1(W2M014),
				.b2(W2M024),
				.b3(W2M104),
				.b4(W2M114),
				.b5(W2M124),
				.b6(W2M204),
				.b7(W2M214),
				.b8(W2M224),
				.c(c2402M)
);

ninexnine_unit ninexnine_unit_6169(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2M005),
				.b1(W2M015),
				.b2(W2M025),
				.b3(W2M105),
				.b4(W2M115),
				.b5(W2M125),
				.b6(W2M205),
				.b7(W2M215),
				.b8(W2M225),
				.c(c2502M)
);

ninexnine_unit ninexnine_unit_6170(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2M006),
				.b1(W2M016),
				.b2(W2M026),
				.b3(W2M106),
				.b4(W2M116),
				.b5(W2M126),
				.b6(W2M206),
				.b7(W2M216),
				.b8(W2M226),
				.c(c2602M)
);

ninexnine_unit ninexnine_unit_6171(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2M007),
				.b1(W2M017),
				.b2(W2M027),
				.b3(W2M107),
				.b4(W2M117),
				.b5(W2M127),
				.b6(W2M207),
				.b7(W2M217),
				.b8(W2M227),
				.c(c2702M)
);

ninexnine_unit ninexnine_unit_6172(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2M008),
				.b1(W2M018),
				.b2(W2M028),
				.b3(W2M108),
				.b4(W2M118),
				.b5(W2M128),
				.b6(W2M208),
				.b7(W2M218),
				.b8(W2M228),
				.c(c2802M)
);

ninexnine_unit ninexnine_unit_6173(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2M009),
				.b1(W2M019),
				.b2(W2M029),
				.b3(W2M109),
				.b4(W2M119),
				.b5(W2M129),
				.b6(W2M209),
				.b7(W2M219),
				.b8(W2M229),
				.c(c2902M)
);

ninexnine_unit ninexnine_unit_6174(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2M00A),
				.b1(W2M01A),
				.b2(W2M02A),
				.b3(W2M10A),
				.b4(W2M11A),
				.b5(W2M12A),
				.b6(W2M20A),
				.b7(W2M21A),
				.b8(W2M22A),
				.c(c2A02M)
);

ninexnine_unit ninexnine_unit_6175(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2M00B),
				.b1(W2M01B),
				.b2(W2M02B),
				.b3(W2M10B),
				.b4(W2M11B),
				.b5(W2M12B),
				.b6(W2M20B),
				.b7(W2M21B),
				.b8(W2M22B),
				.c(c2B02M)
);

ninexnine_unit ninexnine_unit_6176(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2M00C),
				.b1(W2M01C),
				.b2(W2M02C),
				.b3(W2M10C),
				.b4(W2M11C),
				.b5(W2M12C),
				.b6(W2M20C),
				.b7(W2M21C),
				.b8(W2M22C),
				.c(c2C02M)
);

ninexnine_unit ninexnine_unit_6177(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2M00D),
				.b1(W2M01D),
				.b2(W2M02D),
				.b3(W2M10D),
				.b4(W2M11D),
				.b5(W2M12D),
				.b6(W2M20D),
				.b7(W2M21D),
				.b8(W2M22D),
				.c(c2D02M)
);

ninexnine_unit ninexnine_unit_6178(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2M00E),
				.b1(W2M01E),
				.b2(W2M02E),
				.b3(W2M10E),
				.b4(W2M11E),
				.b5(W2M12E),
				.b6(W2M20E),
				.b7(W2M21E),
				.b8(W2M22E),
				.c(c2E02M)
);

ninexnine_unit ninexnine_unit_6179(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2M00F),
				.b1(W2M01F),
				.b2(W2M02F),
				.b3(W2M10F),
				.b4(W2M11F),
				.b5(W2M12F),
				.b6(W2M20F),
				.b7(W2M21F),
				.b8(W2M22F),
				.c(c2F02M)
);

assign C202M=c2002M+c2102M+c2202M+c2302M+c2402M+c2502M+c2602M+c2702M+c2802M+c2902M+c2A02M+c2B02M+c2C02M+c2D02M+c2E02M+c2F02M;
assign A202M=(C202M>=0)?1:0;

assign P302M=A202M;

ninexnine_unit ninexnine_unit_6180(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2M000),
				.b1(W2M010),
				.b2(W2M020),
				.b3(W2M100),
				.b4(W2M110),
				.b5(W2M120),
				.b6(W2M200),
				.b7(W2M210),
				.b8(W2M220),
				.c(c2010M)
);

ninexnine_unit ninexnine_unit_6181(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2M001),
				.b1(W2M011),
				.b2(W2M021),
				.b3(W2M101),
				.b4(W2M111),
				.b5(W2M121),
				.b6(W2M201),
				.b7(W2M211),
				.b8(W2M221),
				.c(c2110M)
);

ninexnine_unit ninexnine_unit_6182(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2M002),
				.b1(W2M012),
				.b2(W2M022),
				.b3(W2M102),
				.b4(W2M112),
				.b5(W2M122),
				.b6(W2M202),
				.b7(W2M212),
				.b8(W2M222),
				.c(c2210M)
);

ninexnine_unit ninexnine_unit_6183(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2M003),
				.b1(W2M013),
				.b2(W2M023),
				.b3(W2M103),
				.b4(W2M113),
				.b5(W2M123),
				.b6(W2M203),
				.b7(W2M213),
				.b8(W2M223),
				.c(c2310M)
);

ninexnine_unit ninexnine_unit_6184(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2M004),
				.b1(W2M014),
				.b2(W2M024),
				.b3(W2M104),
				.b4(W2M114),
				.b5(W2M124),
				.b6(W2M204),
				.b7(W2M214),
				.b8(W2M224),
				.c(c2410M)
);

ninexnine_unit ninexnine_unit_6185(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2M005),
				.b1(W2M015),
				.b2(W2M025),
				.b3(W2M105),
				.b4(W2M115),
				.b5(W2M125),
				.b6(W2M205),
				.b7(W2M215),
				.b8(W2M225),
				.c(c2510M)
);

ninexnine_unit ninexnine_unit_6186(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2M006),
				.b1(W2M016),
				.b2(W2M026),
				.b3(W2M106),
				.b4(W2M116),
				.b5(W2M126),
				.b6(W2M206),
				.b7(W2M216),
				.b8(W2M226),
				.c(c2610M)
);

ninexnine_unit ninexnine_unit_6187(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2M007),
				.b1(W2M017),
				.b2(W2M027),
				.b3(W2M107),
				.b4(W2M117),
				.b5(W2M127),
				.b6(W2M207),
				.b7(W2M217),
				.b8(W2M227),
				.c(c2710M)
);

ninexnine_unit ninexnine_unit_6188(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2M008),
				.b1(W2M018),
				.b2(W2M028),
				.b3(W2M108),
				.b4(W2M118),
				.b5(W2M128),
				.b6(W2M208),
				.b7(W2M218),
				.b8(W2M228),
				.c(c2810M)
);

ninexnine_unit ninexnine_unit_6189(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2M009),
				.b1(W2M019),
				.b2(W2M029),
				.b3(W2M109),
				.b4(W2M119),
				.b5(W2M129),
				.b6(W2M209),
				.b7(W2M219),
				.b8(W2M229),
				.c(c2910M)
);

ninexnine_unit ninexnine_unit_6190(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2M00A),
				.b1(W2M01A),
				.b2(W2M02A),
				.b3(W2M10A),
				.b4(W2M11A),
				.b5(W2M12A),
				.b6(W2M20A),
				.b7(W2M21A),
				.b8(W2M22A),
				.c(c2A10M)
);

ninexnine_unit ninexnine_unit_6191(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2M00B),
				.b1(W2M01B),
				.b2(W2M02B),
				.b3(W2M10B),
				.b4(W2M11B),
				.b5(W2M12B),
				.b6(W2M20B),
				.b7(W2M21B),
				.b8(W2M22B),
				.c(c2B10M)
);

ninexnine_unit ninexnine_unit_6192(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2M00C),
				.b1(W2M01C),
				.b2(W2M02C),
				.b3(W2M10C),
				.b4(W2M11C),
				.b5(W2M12C),
				.b6(W2M20C),
				.b7(W2M21C),
				.b8(W2M22C),
				.c(c2C10M)
);

ninexnine_unit ninexnine_unit_6193(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2M00D),
				.b1(W2M01D),
				.b2(W2M02D),
				.b3(W2M10D),
				.b4(W2M11D),
				.b5(W2M12D),
				.b6(W2M20D),
				.b7(W2M21D),
				.b8(W2M22D),
				.c(c2D10M)
);

ninexnine_unit ninexnine_unit_6194(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2M00E),
				.b1(W2M01E),
				.b2(W2M02E),
				.b3(W2M10E),
				.b4(W2M11E),
				.b5(W2M12E),
				.b6(W2M20E),
				.b7(W2M21E),
				.b8(W2M22E),
				.c(c2E10M)
);

ninexnine_unit ninexnine_unit_6195(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2M00F),
				.b1(W2M01F),
				.b2(W2M02F),
				.b3(W2M10F),
				.b4(W2M11F),
				.b5(W2M12F),
				.b6(W2M20F),
				.b7(W2M21F),
				.b8(W2M22F),
				.c(c2F10M)
);

assign C210M=c2010M+c2110M+c2210M+c2310M+c2410M+c2510M+c2610M+c2710M+c2810M+c2910M+c2A10M+c2B10M+c2C10M+c2D10M+c2E10M+c2F10M;
assign A210M=(C210M>=0)?1:0;

assign P310M=A210M;

ninexnine_unit ninexnine_unit_6196(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2M000),
				.b1(W2M010),
				.b2(W2M020),
				.b3(W2M100),
				.b4(W2M110),
				.b5(W2M120),
				.b6(W2M200),
				.b7(W2M210),
				.b8(W2M220),
				.c(c2011M)
);

ninexnine_unit ninexnine_unit_6197(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2M001),
				.b1(W2M011),
				.b2(W2M021),
				.b3(W2M101),
				.b4(W2M111),
				.b5(W2M121),
				.b6(W2M201),
				.b7(W2M211),
				.b8(W2M221),
				.c(c2111M)
);

ninexnine_unit ninexnine_unit_6198(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2M002),
				.b1(W2M012),
				.b2(W2M022),
				.b3(W2M102),
				.b4(W2M112),
				.b5(W2M122),
				.b6(W2M202),
				.b7(W2M212),
				.b8(W2M222),
				.c(c2211M)
);

ninexnine_unit ninexnine_unit_6199(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2M003),
				.b1(W2M013),
				.b2(W2M023),
				.b3(W2M103),
				.b4(W2M113),
				.b5(W2M123),
				.b6(W2M203),
				.b7(W2M213),
				.b8(W2M223),
				.c(c2311M)
);

ninexnine_unit ninexnine_unit_6200(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2M004),
				.b1(W2M014),
				.b2(W2M024),
				.b3(W2M104),
				.b4(W2M114),
				.b5(W2M124),
				.b6(W2M204),
				.b7(W2M214),
				.b8(W2M224),
				.c(c2411M)
);

ninexnine_unit ninexnine_unit_6201(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2M005),
				.b1(W2M015),
				.b2(W2M025),
				.b3(W2M105),
				.b4(W2M115),
				.b5(W2M125),
				.b6(W2M205),
				.b7(W2M215),
				.b8(W2M225),
				.c(c2511M)
);

ninexnine_unit ninexnine_unit_6202(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2M006),
				.b1(W2M016),
				.b2(W2M026),
				.b3(W2M106),
				.b4(W2M116),
				.b5(W2M126),
				.b6(W2M206),
				.b7(W2M216),
				.b8(W2M226),
				.c(c2611M)
);

ninexnine_unit ninexnine_unit_6203(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2M007),
				.b1(W2M017),
				.b2(W2M027),
				.b3(W2M107),
				.b4(W2M117),
				.b5(W2M127),
				.b6(W2M207),
				.b7(W2M217),
				.b8(W2M227),
				.c(c2711M)
);

ninexnine_unit ninexnine_unit_6204(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2M008),
				.b1(W2M018),
				.b2(W2M028),
				.b3(W2M108),
				.b4(W2M118),
				.b5(W2M128),
				.b6(W2M208),
				.b7(W2M218),
				.b8(W2M228),
				.c(c2811M)
);

ninexnine_unit ninexnine_unit_6205(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2M009),
				.b1(W2M019),
				.b2(W2M029),
				.b3(W2M109),
				.b4(W2M119),
				.b5(W2M129),
				.b6(W2M209),
				.b7(W2M219),
				.b8(W2M229),
				.c(c2911M)
);

ninexnine_unit ninexnine_unit_6206(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2M00A),
				.b1(W2M01A),
				.b2(W2M02A),
				.b3(W2M10A),
				.b4(W2M11A),
				.b5(W2M12A),
				.b6(W2M20A),
				.b7(W2M21A),
				.b8(W2M22A),
				.c(c2A11M)
);

ninexnine_unit ninexnine_unit_6207(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2M00B),
				.b1(W2M01B),
				.b2(W2M02B),
				.b3(W2M10B),
				.b4(W2M11B),
				.b5(W2M12B),
				.b6(W2M20B),
				.b7(W2M21B),
				.b8(W2M22B),
				.c(c2B11M)
);

ninexnine_unit ninexnine_unit_6208(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2M00C),
				.b1(W2M01C),
				.b2(W2M02C),
				.b3(W2M10C),
				.b4(W2M11C),
				.b5(W2M12C),
				.b6(W2M20C),
				.b7(W2M21C),
				.b8(W2M22C),
				.c(c2C11M)
);

ninexnine_unit ninexnine_unit_6209(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2M00D),
				.b1(W2M01D),
				.b2(W2M02D),
				.b3(W2M10D),
				.b4(W2M11D),
				.b5(W2M12D),
				.b6(W2M20D),
				.b7(W2M21D),
				.b8(W2M22D),
				.c(c2D11M)
);

ninexnine_unit ninexnine_unit_6210(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2M00E),
				.b1(W2M01E),
				.b2(W2M02E),
				.b3(W2M10E),
				.b4(W2M11E),
				.b5(W2M12E),
				.b6(W2M20E),
				.b7(W2M21E),
				.b8(W2M22E),
				.c(c2E11M)
);

ninexnine_unit ninexnine_unit_6211(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2M00F),
				.b1(W2M01F),
				.b2(W2M02F),
				.b3(W2M10F),
				.b4(W2M11F),
				.b5(W2M12F),
				.b6(W2M20F),
				.b7(W2M21F),
				.b8(W2M22F),
				.c(c2F11M)
);

assign C211M=c2011M+c2111M+c2211M+c2311M+c2411M+c2511M+c2611M+c2711M+c2811M+c2911M+c2A11M+c2B11M+c2C11M+c2D11M+c2E11M+c2F11M;
assign A211M=(C211M>=0)?1:0;

assign P311M=A211M;

ninexnine_unit ninexnine_unit_6212(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2M000),
				.b1(W2M010),
				.b2(W2M020),
				.b3(W2M100),
				.b4(W2M110),
				.b5(W2M120),
				.b6(W2M200),
				.b7(W2M210),
				.b8(W2M220),
				.c(c2012M)
);

ninexnine_unit ninexnine_unit_6213(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2M001),
				.b1(W2M011),
				.b2(W2M021),
				.b3(W2M101),
				.b4(W2M111),
				.b5(W2M121),
				.b6(W2M201),
				.b7(W2M211),
				.b8(W2M221),
				.c(c2112M)
);

ninexnine_unit ninexnine_unit_6214(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2M002),
				.b1(W2M012),
				.b2(W2M022),
				.b3(W2M102),
				.b4(W2M112),
				.b5(W2M122),
				.b6(W2M202),
				.b7(W2M212),
				.b8(W2M222),
				.c(c2212M)
);

ninexnine_unit ninexnine_unit_6215(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2M003),
				.b1(W2M013),
				.b2(W2M023),
				.b3(W2M103),
				.b4(W2M113),
				.b5(W2M123),
				.b6(W2M203),
				.b7(W2M213),
				.b8(W2M223),
				.c(c2312M)
);

ninexnine_unit ninexnine_unit_6216(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2M004),
				.b1(W2M014),
				.b2(W2M024),
				.b3(W2M104),
				.b4(W2M114),
				.b5(W2M124),
				.b6(W2M204),
				.b7(W2M214),
				.b8(W2M224),
				.c(c2412M)
);

ninexnine_unit ninexnine_unit_6217(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2M005),
				.b1(W2M015),
				.b2(W2M025),
				.b3(W2M105),
				.b4(W2M115),
				.b5(W2M125),
				.b6(W2M205),
				.b7(W2M215),
				.b8(W2M225),
				.c(c2512M)
);

ninexnine_unit ninexnine_unit_6218(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2M006),
				.b1(W2M016),
				.b2(W2M026),
				.b3(W2M106),
				.b4(W2M116),
				.b5(W2M126),
				.b6(W2M206),
				.b7(W2M216),
				.b8(W2M226),
				.c(c2612M)
);

ninexnine_unit ninexnine_unit_6219(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2M007),
				.b1(W2M017),
				.b2(W2M027),
				.b3(W2M107),
				.b4(W2M117),
				.b5(W2M127),
				.b6(W2M207),
				.b7(W2M217),
				.b8(W2M227),
				.c(c2712M)
);

ninexnine_unit ninexnine_unit_6220(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2M008),
				.b1(W2M018),
				.b2(W2M028),
				.b3(W2M108),
				.b4(W2M118),
				.b5(W2M128),
				.b6(W2M208),
				.b7(W2M218),
				.b8(W2M228),
				.c(c2812M)
);

ninexnine_unit ninexnine_unit_6221(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2M009),
				.b1(W2M019),
				.b2(W2M029),
				.b3(W2M109),
				.b4(W2M119),
				.b5(W2M129),
				.b6(W2M209),
				.b7(W2M219),
				.b8(W2M229),
				.c(c2912M)
);

ninexnine_unit ninexnine_unit_6222(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2M00A),
				.b1(W2M01A),
				.b2(W2M02A),
				.b3(W2M10A),
				.b4(W2M11A),
				.b5(W2M12A),
				.b6(W2M20A),
				.b7(W2M21A),
				.b8(W2M22A),
				.c(c2A12M)
);

ninexnine_unit ninexnine_unit_6223(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2M00B),
				.b1(W2M01B),
				.b2(W2M02B),
				.b3(W2M10B),
				.b4(W2M11B),
				.b5(W2M12B),
				.b6(W2M20B),
				.b7(W2M21B),
				.b8(W2M22B),
				.c(c2B12M)
);

ninexnine_unit ninexnine_unit_6224(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2M00C),
				.b1(W2M01C),
				.b2(W2M02C),
				.b3(W2M10C),
				.b4(W2M11C),
				.b5(W2M12C),
				.b6(W2M20C),
				.b7(W2M21C),
				.b8(W2M22C),
				.c(c2C12M)
);

ninexnine_unit ninexnine_unit_6225(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2M00D),
				.b1(W2M01D),
				.b2(W2M02D),
				.b3(W2M10D),
				.b4(W2M11D),
				.b5(W2M12D),
				.b6(W2M20D),
				.b7(W2M21D),
				.b8(W2M22D),
				.c(c2D12M)
);

ninexnine_unit ninexnine_unit_6226(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2M00E),
				.b1(W2M01E),
				.b2(W2M02E),
				.b3(W2M10E),
				.b4(W2M11E),
				.b5(W2M12E),
				.b6(W2M20E),
				.b7(W2M21E),
				.b8(W2M22E),
				.c(c2E12M)
);

ninexnine_unit ninexnine_unit_6227(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2M00F),
				.b1(W2M01F),
				.b2(W2M02F),
				.b3(W2M10F),
				.b4(W2M11F),
				.b5(W2M12F),
				.b6(W2M20F),
				.b7(W2M21F),
				.b8(W2M22F),
				.c(c2F12M)
);

assign C212M=c2012M+c2112M+c2212M+c2312M+c2412M+c2512M+c2612M+c2712M+c2812M+c2912M+c2A12M+c2B12M+c2C12M+c2D12M+c2E12M+c2F12M;
assign A212M=(C212M>=0)?1:0;

assign P312M=A212M;

ninexnine_unit ninexnine_unit_6228(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2M000),
				.b1(W2M010),
				.b2(W2M020),
				.b3(W2M100),
				.b4(W2M110),
				.b5(W2M120),
				.b6(W2M200),
				.b7(W2M210),
				.b8(W2M220),
				.c(c2020M)
);

ninexnine_unit ninexnine_unit_6229(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2M001),
				.b1(W2M011),
				.b2(W2M021),
				.b3(W2M101),
				.b4(W2M111),
				.b5(W2M121),
				.b6(W2M201),
				.b7(W2M211),
				.b8(W2M221),
				.c(c2120M)
);

ninexnine_unit ninexnine_unit_6230(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2M002),
				.b1(W2M012),
				.b2(W2M022),
				.b3(W2M102),
				.b4(W2M112),
				.b5(W2M122),
				.b6(W2M202),
				.b7(W2M212),
				.b8(W2M222),
				.c(c2220M)
);

ninexnine_unit ninexnine_unit_6231(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2M003),
				.b1(W2M013),
				.b2(W2M023),
				.b3(W2M103),
				.b4(W2M113),
				.b5(W2M123),
				.b6(W2M203),
				.b7(W2M213),
				.b8(W2M223),
				.c(c2320M)
);

ninexnine_unit ninexnine_unit_6232(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2M004),
				.b1(W2M014),
				.b2(W2M024),
				.b3(W2M104),
				.b4(W2M114),
				.b5(W2M124),
				.b6(W2M204),
				.b7(W2M214),
				.b8(W2M224),
				.c(c2420M)
);

ninexnine_unit ninexnine_unit_6233(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2M005),
				.b1(W2M015),
				.b2(W2M025),
				.b3(W2M105),
				.b4(W2M115),
				.b5(W2M125),
				.b6(W2M205),
				.b7(W2M215),
				.b8(W2M225),
				.c(c2520M)
);

ninexnine_unit ninexnine_unit_6234(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2M006),
				.b1(W2M016),
				.b2(W2M026),
				.b3(W2M106),
				.b4(W2M116),
				.b5(W2M126),
				.b6(W2M206),
				.b7(W2M216),
				.b8(W2M226),
				.c(c2620M)
);

ninexnine_unit ninexnine_unit_6235(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2M007),
				.b1(W2M017),
				.b2(W2M027),
				.b3(W2M107),
				.b4(W2M117),
				.b5(W2M127),
				.b6(W2M207),
				.b7(W2M217),
				.b8(W2M227),
				.c(c2720M)
);

ninexnine_unit ninexnine_unit_6236(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2M008),
				.b1(W2M018),
				.b2(W2M028),
				.b3(W2M108),
				.b4(W2M118),
				.b5(W2M128),
				.b6(W2M208),
				.b7(W2M218),
				.b8(W2M228),
				.c(c2820M)
);

ninexnine_unit ninexnine_unit_6237(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2M009),
				.b1(W2M019),
				.b2(W2M029),
				.b3(W2M109),
				.b4(W2M119),
				.b5(W2M129),
				.b6(W2M209),
				.b7(W2M219),
				.b8(W2M229),
				.c(c2920M)
);

ninexnine_unit ninexnine_unit_6238(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2M00A),
				.b1(W2M01A),
				.b2(W2M02A),
				.b3(W2M10A),
				.b4(W2M11A),
				.b5(W2M12A),
				.b6(W2M20A),
				.b7(W2M21A),
				.b8(W2M22A),
				.c(c2A20M)
);

ninexnine_unit ninexnine_unit_6239(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2M00B),
				.b1(W2M01B),
				.b2(W2M02B),
				.b3(W2M10B),
				.b4(W2M11B),
				.b5(W2M12B),
				.b6(W2M20B),
				.b7(W2M21B),
				.b8(W2M22B),
				.c(c2B20M)
);

ninexnine_unit ninexnine_unit_6240(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2M00C),
				.b1(W2M01C),
				.b2(W2M02C),
				.b3(W2M10C),
				.b4(W2M11C),
				.b5(W2M12C),
				.b6(W2M20C),
				.b7(W2M21C),
				.b8(W2M22C),
				.c(c2C20M)
);

ninexnine_unit ninexnine_unit_6241(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2M00D),
				.b1(W2M01D),
				.b2(W2M02D),
				.b3(W2M10D),
				.b4(W2M11D),
				.b5(W2M12D),
				.b6(W2M20D),
				.b7(W2M21D),
				.b8(W2M22D),
				.c(c2D20M)
);

ninexnine_unit ninexnine_unit_6242(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2M00E),
				.b1(W2M01E),
				.b2(W2M02E),
				.b3(W2M10E),
				.b4(W2M11E),
				.b5(W2M12E),
				.b6(W2M20E),
				.b7(W2M21E),
				.b8(W2M22E),
				.c(c2E20M)
);

ninexnine_unit ninexnine_unit_6243(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2M00F),
				.b1(W2M01F),
				.b2(W2M02F),
				.b3(W2M10F),
				.b4(W2M11F),
				.b5(W2M12F),
				.b6(W2M20F),
				.b7(W2M21F),
				.b8(W2M22F),
				.c(c2F20M)
);

assign C220M=c2020M+c2120M+c2220M+c2320M+c2420M+c2520M+c2620M+c2720M+c2820M+c2920M+c2A20M+c2B20M+c2C20M+c2D20M+c2E20M+c2F20M;
assign A220M=(C220M>=0)?1:0;

assign P320M=A220M;

ninexnine_unit ninexnine_unit_6244(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2M000),
				.b1(W2M010),
				.b2(W2M020),
				.b3(W2M100),
				.b4(W2M110),
				.b5(W2M120),
				.b6(W2M200),
				.b7(W2M210),
				.b8(W2M220),
				.c(c2021M)
);

ninexnine_unit ninexnine_unit_6245(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2M001),
				.b1(W2M011),
				.b2(W2M021),
				.b3(W2M101),
				.b4(W2M111),
				.b5(W2M121),
				.b6(W2M201),
				.b7(W2M211),
				.b8(W2M221),
				.c(c2121M)
);

ninexnine_unit ninexnine_unit_6246(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2M002),
				.b1(W2M012),
				.b2(W2M022),
				.b3(W2M102),
				.b4(W2M112),
				.b5(W2M122),
				.b6(W2M202),
				.b7(W2M212),
				.b8(W2M222),
				.c(c2221M)
);

ninexnine_unit ninexnine_unit_6247(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2M003),
				.b1(W2M013),
				.b2(W2M023),
				.b3(W2M103),
				.b4(W2M113),
				.b5(W2M123),
				.b6(W2M203),
				.b7(W2M213),
				.b8(W2M223),
				.c(c2321M)
);

ninexnine_unit ninexnine_unit_6248(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2M004),
				.b1(W2M014),
				.b2(W2M024),
				.b3(W2M104),
				.b4(W2M114),
				.b5(W2M124),
				.b6(W2M204),
				.b7(W2M214),
				.b8(W2M224),
				.c(c2421M)
);

ninexnine_unit ninexnine_unit_6249(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2M005),
				.b1(W2M015),
				.b2(W2M025),
				.b3(W2M105),
				.b4(W2M115),
				.b5(W2M125),
				.b6(W2M205),
				.b7(W2M215),
				.b8(W2M225),
				.c(c2521M)
);

ninexnine_unit ninexnine_unit_6250(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2M006),
				.b1(W2M016),
				.b2(W2M026),
				.b3(W2M106),
				.b4(W2M116),
				.b5(W2M126),
				.b6(W2M206),
				.b7(W2M216),
				.b8(W2M226),
				.c(c2621M)
);

ninexnine_unit ninexnine_unit_6251(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2M007),
				.b1(W2M017),
				.b2(W2M027),
				.b3(W2M107),
				.b4(W2M117),
				.b5(W2M127),
				.b6(W2M207),
				.b7(W2M217),
				.b8(W2M227),
				.c(c2721M)
);

ninexnine_unit ninexnine_unit_6252(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2M008),
				.b1(W2M018),
				.b2(W2M028),
				.b3(W2M108),
				.b4(W2M118),
				.b5(W2M128),
				.b6(W2M208),
				.b7(W2M218),
				.b8(W2M228),
				.c(c2821M)
);

ninexnine_unit ninexnine_unit_6253(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2M009),
				.b1(W2M019),
				.b2(W2M029),
				.b3(W2M109),
				.b4(W2M119),
				.b5(W2M129),
				.b6(W2M209),
				.b7(W2M219),
				.b8(W2M229),
				.c(c2921M)
);

ninexnine_unit ninexnine_unit_6254(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2M00A),
				.b1(W2M01A),
				.b2(W2M02A),
				.b3(W2M10A),
				.b4(W2M11A),
				.b5(W2M12A),
				.b6(W2M20A),
				.b7(W2M21A),
				.b8(W2M22A),
				.c(c2A21M)
);

ninexnine_unit ninexnine_unit_6255(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2M00B),
				.b1(W2M01B),
				.b2(W2M02B),
				.b3(W2M10B),
				.b4(W2M11B),
				.b5(W2M12B),
				.b6(W2M20B),
				.b7(W2M21B),
				.b8(W2M22B),
				.c(c2B21M)
);

ninexnine_unit ninexnine_unit_6256(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2M00C),
				.b1(W2M01C),
				.b2(W2M02C),
				.b3(W2M10C),
				.b4(W2M11C),
				.b5(W2M12C),
				.b6(W2M20C),
				.b7(W2M21C),
				.b8(W2M22C),
				.c(c2C21M)
);

ninexnine_unit ninexnine_unit_6257(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2M00D),
				.b1(W2M01D),
				.b2(W2M02D),
				.b3(W2M10D),
				.b4(W2M11D),
				.b5(W2M12D),
				.b6(W2M20D),
				.b7(W2M21D),
				.b8(W2M22D),
				.c(c2D21M)
);

ninexnine_unit ninexnine_unit_6258(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2M00E),
				.b1(W2M01E),
				.b2(W2M02E),
				.b3(W2M10E),
				.b4(W2M11E),
				.b5(W2M12E),
				.b6(W2M20E),
				.b7(W2M21E),
				.b8(W2M22E),
				.c(c2E21M)
);

ninexnine_unit ninexnine_unit_6259(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2M00F),
				.b1(W2M01F),
				.b2(W2M02F),
				.b3(W2M10F),
				.b4(W2M11F),
				.b5(W2M12F),
				.b6(W2M20F),
				.b7(W2M21F),
				.b8(W2M22F),
				.c(c2F21M)
);

assign C221M=c2021M+c2121M+c2221M+c2321M+c2421M+c2521M+c2621M+c2721M+c2821M+c2921M+c2A21M+c2B21M+c2C21M+c2D21M+c2E21M+c2F21M;
assign A221M=(C221M>=0)?1:0;

assign P321M=A221M;

ninexnine_unit ninexnine_unit_6260(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2M000),
				.b1(W2M010),
				.b2(W2M020),
				.b3(W2M100),
				.b4(W2M110),
				.b5(W2M120),
				.b6(W2M200),
				.b7(W2M210),
				.b8(W2M220),
				.c(c2022M)
);

ninexnine_unit ninexnine_unit_6261(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2M001),
				.b1(W2M011),
				.b2(W2M021),
				.b3(W2M101),
				.b4(W2M111),
				.b5(W2M121),
				.b6(W2M201),
				.b7(W2M211),
				.b8(W2M221),
				.c(c2122M)
);

ninexnine_unit ninexnine_unit_6262(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2M002),
				.b1(W2M012),
				.b2(W2M022),
				.b3(W2M102),
				.b4(W2M112),
				.b5(W2M122),
				.b6(W2M202),
				.b7(W2M212),
				.b8(W2M222),
				.c(c2222M)
);

ninexnine_unit ninexnine_unit_6263(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2M003),
				.b1(W2M013),
				.b2(W2M023),
				.b3(W2M103),
				.b4(W2M113),
				.b5(W2M123),
				.b6(W2M203),
				.b7(W2M213),
				.b8(W2M223),
				.c(c2322M)
);

ninexnine_unit ninexnine_unit_6264(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2M004),
				.b1(W2M014),
				.b2(W2M024),
				.b3(W2M104),
				.b4(W2M114),
				.b5(W2M124),
				.b6(W2M204),
				.b7(W2M214),
				.b8(W2M224),
				.c(c2422M)
);

ninexnine_unit ninexnine_unit_6265(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2M005),
				.b1(W2M015),
				.b2(W2M025),
				.b3(W2M105),
				.b4(W2M115),
				.b5(W2M125),
				.b6(W2M205),
				.b7(W2M215),
				.b8(W2M225),
				.c(c2522M)
);

ninexnine_unit ninexnine_unit_6266(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2M006),
				.b1(W2M016),
				.b2(W2M026),
				.b3(W2M106),
				.b4(W2M116),
				.b5(W2M126),
				.b6(W2M206),
				.b7(W2M216),
				.b8(W2M226),
				.c(c2622M)
);

ninexnine_unit ninexnine_unit_6267(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2M007),
				.b1(W2M017),
				.b2(W2M027),
				.b3(W2M107),
				.b4(W2M117),
				.b5(W2M127),
				.b6(W2M207),
				.b7(W2M217),
				.b8(W2M227),
				.c(c2722M)
);

ninexnine_unit ninexnine_unit_6268(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2M008),
				.b1(W2M018),
				.b2(W2M028),
				.b3(W2M108),
				.b4(W2M118),
				.b5(W2M128),
				.b6(W2M208),
				.b7(W2M218),
				.b8(W2M228),
				.c(c2822M)
);

ninexnine_unit ninexnine_unit_6269(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2M009),
				.b1(W2M019),
				.b2(W2M029),
				.b3(W2M109),
				.b4(W2M119),
				.b5(W2M129),
				.b6(W2M209),
				.b7(W2M219),
				.b8(W2M229),
				.c(c2922M)
);

ninexnine_unit ninexnine_unit_6270(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2M00A),
				.b1(W2M01A),
				.b2(W2M02A),
				.b3(W2M10A),
				.b4(W2M11A),
				.b5(W2M12A),
				.b6(W2M20A),
				.b7(W2M21A),
				.b8(W2M22A),
				.c(c2A22M)
);

ninexnine_unit ninexnine_unit_6271(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2M00B),
				.b1(W2M01B),
				.b2(W2M02B),
				.b3(W2M10B),
				.b4(W2M11B),
				.b5(W2M12B),
				.b6(W2M20B),
				.b7(W2M21B),
				.b8(W2M22B),
				.c(c2B22M)
);

ninexnine_unit ninexnine_unit_6272(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2M00C),
				.b1(W2M01C),
				.b2(W2M02C),
				.b3(W2M10C),
				.b4(W2M11C),
				.b5(W2M12C),
				.b6(W2M20C),
				.b7(W2M21C),
				.b8(W2M22C),
				.c(c2C22M)
);

ninexnine_unit ninexnine_unit_6273(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2M00D),
				.b1(W2M01D),
				.b2(W2M02D),
				.b3(W2M10D),
				.b4(W2M11D),
				.b5(W2M12D),
				.b6(W2M20D),
				.b7(W2M21D),
				.b8(W2M22D),
				.c(c2D22M)
);

ninexnine_unit ninexnine_unit_6274(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2M00E),
				.b1(W2M01E),
				.b2(W2M02E),
				.b3(W2M10E),
				.b4(W2M11E),
				.b5(W2M12E),
				.b6(W2M20E),
				.b7(W2M21E),
				.b8(W2M22E),
				.c(c2E22M)
);

ninexnine_unit ninexnine_unit_6275(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2M00F),
				.b1(W2M01F),
				.b2(W2M02F),
				.b3(W2M10F),
				.b4(W2M11F),
				.b5(W2M12F),
				.b6(W2M20F),
				.b7(W2M21F),
				.b8(W2M22F),
				.c(c2F22M)
);

assign C222M=c2022M+c2122M+c2222M+c2322M+c2422M+c2522M+c2622M+c2722M+c2822M+c2922M+c2A22M+c2B22M+c2C22M+c2D22M+c2E22M+c2F22M;
assign A222M=(C222M>=0)?1:0;

assign P322M=A222M;

ninexnine_unit ninexnine_unit_6276(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2N000),
				.b1(W2N010),
				.b2(W2N020),
				.b3(W2N100),
				.b4(W2N110),
				.b5(W2N120),
				.b6(W2N200),
				.b7(W2N210),
				.b8(W2N220),
				.c(c2000N)
);

ninexnine_unit ninexnine_unit_6277(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2N001),
				.b1(W2N011),
				.b2(W2N021),
				.b3(W2N101),
				.b4(W2N111),
				.b5(W2N121),
				.b6(W2N201),
				.b7(W2N211),
				.b8(W2N221),
				.c(c2100N)
);

ninexnine_unit ninexnine_unit_6278(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2N002),
				.b1(W2N012),
				.b2(W2N022),
				.b3(W2N102),
				.b4(W2N112),
				.b5(W2N122),
				.b6(W2N202),
				.b7(W2N212),
				.b8(W2N222),
				.c(c2200N)
);

ninexnine_unit ninexnine_unit_6279(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2N003),
				.b1(W2N013),
				.b2(W2N023),
				.b3(W2N103),
				.b4(W2N113),
				.b5(W2N123),
				.b6(W2N203),
				.b7(W2N213),
				.b8(W2N223),
				.c(c2300N)
);

ninexnine_unit ninexnine_unit_6280(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2N004),
				.b1(W2N014),
				.b2(W2N024),
				.b3(W2N104),
				.b4(W2N114),
				.b5(W2N124),
				.b6(W2N204),
				.b7(W2N214),
				.b8(W2N224),
				.c(c2400N)
);

ninexnine_unit ninexnine_unit_6281(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2N005),
				.b1(W2N015),
				.b2(W2N025),
				.b3(W2N105),
				.b4(W2N115),
				.b5(W2N125),
				.b6(W2N205),
				.b7(W2N215),
				.b8(W2N225),
				.c(c2500N)
);

ninexnine_unit ninexnine_unit_6282(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2N006),
				.b1(W2N016),
				.b2(W2N026),
				.b3(W2N106),
				.b4(W2N116),
				.b5(W2N126),
				.b6(W2N206),
				.b7(W2N216),
				.b8(W2N226),
				.c(c2600N)
);

ninexnine_unit ninexnine_unit_6283(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2N007),
				.b1(W2N017),
				.b2(W2N027),
				.b3(W2N107),
				.b4(W2N117),
				.b5(W2N127),
				.b6(W2N207),
				.b7(W2N217),
				.b8(W2N227),
				.c(c2700N)
);

ninexnine_unit ninexnine_unit_6284(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2N008),
				.b1(W2N018),
				.b2(W2N028),
				.b3(W2N108),
				.b4(W2N118),
				.b5(W2N128),
				.b6(W2N208),
				.b7(W2N218),
				.b8(W2N228),
				.c(c2800N)
);

ninexnine_unit ninexnine_unit_6285(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2N009),
				.b1(W2N019),
				.b2(W2N029),
				.b3(W2N109),
				.b4(W2N119),
				.b5(W2N129),
				.b6(W2N209),
				.b7(W2N219),
				.b8(W2N229),
				.c(c2900N)
);

ninexnine_unit ninexnine_unit_6286(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2N00A),
				.b1(W2N01A),
				.b2(W2N02A),
				.b3(W2N10A),
				.b4(W2N11A),
				.b5(W2N12A),
				.b6(W2N20A),
				.b7(W2N21A),
				.b8(W2N22A),
				.c(c2A00N)
);

ninexnine_unit ninexnine_unit_6287(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2N00B),
				.b1(W2N01B),
				.b2(W2N02B),
				.b3(W2N10B),
				.b4(W2N11B),
				.b5(W2N12B),
				.b6(W2N20B),
				.b7(W2N21B),
				.b8(W2N22B),
				.c(c2B00N)
);

ninexnine_unit ninexnine_unit_6288(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2N00C),
				.b1(W2N01C),
				.b2(W2N02C),
				.b3(W2N10C),
				.b4(W2N11C),
				.b5(W2N12C),
				.b6(W2N20C),
				.b7(W2N21C),
				.b8(W2N22C),
				.c(c2C00N)
);

ninexnine_unit ninexnine_unit_6289(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2N00D),
				.b1(W2N01D),
				.b2(W2N02D),
				.b3(W2N10D),
				.b4(W2N11D),
				.b5(W2N12D),
				.b6(W2N20D),
				.b7(W2N21D),
				.b8(W2N22D),
				.c(c2D00N)
);

ninexnine_unit ninexnine_unit_6290(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2N00E),
				.b1(W2N01E),
				.b2(W2N02E),
				.b3(W2N10E),
				.b4(W2N11E),
				.b5(W2N12E),
				.b6(W2N20E),
				.b7(W2N21E),
				.b8(W2N22E),
				.c(c2E00N)
);

ninexnine_unit ninexnine_unit_6291(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2N00F),
				.b1(W2N01F),
				.b2(W2N02F),
				.b3(W2N10F),
				.b4(W2N11F),
				.b5(W2N12F),
				.b6(W2N20F),
				.b7(W2N21F),
				.b8(W2N22F),
				.c(c2F00N)
);

assign C200N=c2000N+c2100N+c2200N+c2300N+c2400N+c2500N+c2600N+c2700N+c2800N+c2900N+c2A00N+c2B00N+c2C00N+c2D00N+c2E00N+c2F00N;
assign A200N=(C200N>=0)?1:0;

assign P300N=A200N;

ninexnine_unit ninexnine_unit_6292(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2N000),
				.b1(W2N010),
				.b2(W2N020),
				.b3(W2N100),
				.b4(W2N110),
				.b5(W2N120),
				.b6(W2N200),
				.b7(W2N210),
				.b8(W2N220),
				.c(c2001N)
);

ninexnine_unit ninexnine_unit_6293(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2N001),
				.b1(W2N011),
				.b2(W2N021),
				.b3(W2N101),
				.b4(W2N111),
				.b5(W2N121),
				.b6(W2N201),
				.b7(W2N211),
				.b8(W2N221),
				.c(c2101N)
);

ninexnine_unit ninexnine_unit_6294(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2N002),
				.b1(W2N012),
				.b2(W2N022),
				.b3(W2N102),
				.b4(W2N112),
				.b5(W2N122),
				.b6(W2N202),
				.b7(W2N212),
				.b8(W2N222),
				.c(c2201N)
);

ninexnine_unit ninexnine_unit_6295(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2N003),
				.b1(W2N013),
				.b2(W2N023),
				.b3(W2N103),
				.b4(W2N113),
				.b5(W2N123),
				.b6(W2N203),
				.b7(W2N213),
				.b8(W2N223),
				.c(c2301N)
);

ninexnine_unit ninexnine_unit_6296(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2N004),
				.b1(W2N014),
				.b2(W2N024),
				.b3(W2N104),
				.b4(W2N114),
				.b5(W2N124),
				.b6(W2N204),
				.b7(W2N214),
				.b8(W2N224),
				.c(c2401N)
);

ninexnine_unit ninexnine_unit_6297(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2N005),
				.b1(W2N015),
				.b2(W2N025),
				.b3(W2N105),
				.b4(W2N115),
				.b5(W2N125),
				.b6(W2N205),
				.b7(W2N215),
				.b8(W2N225),
				.c(c2501N)
);

ninexnine_unit ninexnine_unit_6298(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2N006),
				.b1(W2N016),
				.b2(W2N026),
				.b3(W2N106),
				.b4(W2N116),
				.b5(W2N126),
				.b6(W2N206),
				.b7(W2N216),
				.b8(W2N226),
				.c(c2601N)
);

ninexnine_unit ninexnine_unit_6299(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2N007),
				.b1(W2N017),
				.b2(W2N027),
				.b3(W2N107),
				.b4(W2N117),
				.b5(W2N127),
				.b6(W2N207),
				.b7(W2N217),
				.b8(W2N227),
				.c(c2701N)
);

ninexnine_unit ninexnine_unit_6300(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2N008),
				.b1(W2N018),
				.b2(W2N028),
				.b3(W2N108),
				.b4(W2N118),
				.b5(W2N128),
				.b6(W2N208),
				.b7(W2N218),
				.b8(W2N228),
				.c(c2801N)
);

ninexnine_unit ninexnine_unit_6301(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2N009),
				.b1(W2N019),
				.b2(W2N029),
				.b3(W2N109),
				.b4(W2N119),
				.b5(W2N129),
				.b6(W2N209),
				.b7(W2N219),
				.b8(W2N229),
				.c(c2901N)
);

ninexnine_unit ninexnine_unit_6302(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2N00A),
				.b1(W2N01A),
				.b2(W2N02A),
				.b3(W2N10A),
				.b4(W2N11A),
				.b5(W2N12A),
				.b6(W2N20A),
				.b7(W2N21A),
				.b8(W2N22A),
				.c(c2A01N)
);

ninexnine_unit ninexnine_unit_6303(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2N00B),
				.b1(W2N01B),
				.b2(W2N02B),
				.b3(W2N10B),
				.b4(W2N11B),
				.b5(W2N12B),
				.b6(W2N20B),
				.b7(W2N21B),
				.b8(W2N22B),
				.c(c2B01N)
);

ninexnine_unit ninexnine_unit_6304(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2N00C),
				.b1(W2N01C),
				.b2(W2N02C),
				.b3(W2N10C),
				.b4(W2N11C),
				.b5(W2N12C),
				.b6(W2N20C),
				.b7(W2N21C),
				.b8(W2N22C),
				.c(c2C01N)
);

ninexnine_unit ninexnine_unit_6305(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2N00D),
				.b1(W2N01D),
				.b2(W2N02D),
				.b3(W2N10D),
				.b4(W2N11D),
				.b5(W2N12D),
				.b6(W2N20D),
				.b7(W2N21D),
				.b8(W2N22D),
				.c(c2D01N)
);

ninexnine_unit ninexnine_unit_6306(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2N00E),
				.b1(W2N01E),
				.b2(W2N02E),
				.b3(W2N10E),
				.b4(W2N11E),
				.b5(W2N12E),
				.b6(W2N20E),
				.b7(W2N21E),
				.b8(W2N22E),
				.c(c2E01N)
);

ninexnine_unit ninexnine_unit_6307(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2N00F),
				.b1(W2N01F),
				.b2(W2N02F),
				.b3(W2N10F),
				.b4(W2N11F),
				.b5(W2N12F),
				.b6(W2N20F),
				.b7(W2N21F),
				.b8(W2N22F),
				.c(c2F01N)
);

assign C201N=c2001N+c2101N+c2201N+c2301N+c2401N+c2501N+c2601N+c2701N+c2801N+c2901N+c2A01N+c2B01N+c2C01N+c2D01N+c2E01N+c2F01N;
assign A201N=(C201N>=0)?1:0;

assign P301N=A201N;

ninexnine_unit ninexnine_unit_6308(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2N000),
				.b1(W2N010),
				.b2(W2N020),
				.b3(W2N100),
				.b4(W2N110),
				.b5(W2N120),
				.b6(W2N200),
				.b7(W2N210),
				.b8(W2N220),
				.c(c2002N)
);

ninexnine_unit ninexnine_unit_6309(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2N001),
				.b1(W2N011),
				.b2(W2N021),
				.b3(W2N101),
				.b4(W2N111),
				.b5(W2N121),
				.b6(W2N201),
				.b7(W2N211),
				.b8(W2N221),
				.c(c2102N)
);

ninexnine_unit ninexnine_unit_6310(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2N002),
				.b1(W2N012),
				.b2(W2N022),
				.b3(W2N102),
				.b4(W2N112),
				.b5(W2N122),
				.b6(W2N202),
				.b7(W2N212),
				.b8(W2N222),
				.c(c2202N)
);

ninexnine_unit ninexnine_unit_6311(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2N003),
				.b1(W2N013),
				.b2(W2N023),
				.b3(W2N103),
				.b4(W2N113),
				.b5(W2N123),
				.b6(W2N203),
				.b7(W2N213),
				.b8(W2N223),
				.c(c2302N)
);

ninexnine_unit ninexnine_unit_6312(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2N004),
				.b1(W2N014),
				.b2(W2N024),
				.b3(W2N104),
				.b4(W2N114),
				.b5(W2N124),
				.b6(W2N204),
				.b7(W2N214),
				.b8(W2N224),
				.c(c2402N)
);

ninexnine_unit ninexnine_unit_6313(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2N005),
				.b1(W2N015),
				.b2(W2N025),
				.b3(W2N105),
				.b4(W2N115),
				.b5(W2N125),
				.b6(W2N205),
				.b7(W2N215),
				.b8(W2N225),
				.c(c2502N)
);

ninexnine_unit ninexnine_unit_6314(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2N006),
				.b1(W2N016),
				.b2(W2N026),
				.b3(W2N106),
				.b4(W2N116),
				.b5(W2N126),
				.b6(W2N206),
				.b7(W2N216),
				.b8(W2N226),
				.c(c2602N)
);

ninexnine_unit ninexnine_unit_6315(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2N007),
				.b1(W2N017),
				.b2(W2N027),
				.b3(W2N107),
				.b4(W2N117),
				.b5(W2N127),
				.b6(W2N207),
				.b7(W2N217),
				.b8(W2N227),
				.c(c2702N)
);

ninexnine_unit ninexnine_unit_6316(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2N008),
				.b1(W2N018),
				.b2(W2N028),
				.b3(W2N108),
				.b4(W2N118),
				.b5(W2N128),
				.b6(W2N208),
				.b7(W2N218),
				.b8(W2N228),
				.c(c2802N)
);

ninexnine_unit ninexnine_unit_6317(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2N009),
				.b1(W2N019),
				.b2(W2N029),
				.b3(W2N109),
				.b4(W2N119),
				.b5(W2N129),
				.b6(W2N209),
				.b7(W2N219),
				.b8(W2N229),
				.c(c2902N)
);

ninexnine_unit ninexnine_unit_6318(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2N00A),
				.b1(W2N01A),
				.b2(W2N02A),
				.b3(W2N10A),
				.b4(W2N11A),
				.b5(W2N12A),
				.b6(W2N20A),
				.b7(W2N21A),
				.b8(W2N22A),
				.c(c2A02N)
);

ninexnine_unit ninexnine_unit_6319(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2N00B),
				.b1(W2N01B),
				.b2(W2N02B),
				.b3(W2N10B),
				.b4(W2N11B),
				.b5(W2N12B),
				.b6(W2N20B),
				.b7(W2N21B),
				.b8(W2N22B),
				.c(c2B02N)
);

ninexnine_unit ninexnine_unit_6320(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2N00C),
				.b1(W2N01C),
				.b2(W2N02C),
				.b3(W2N10C),
				.b4(W2N11C),
				.b5(W2N12C),
				.b6(W2N20C),
				.b7(W2N21C),
				.b8(W2N22C),
				.c(c2C02N)
);

ninexnine_unit ninexnine_unit_6321(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2N00D),
				.b1(W2N01D),
				.b2(W2N02D),
				.b3(W2N10D),
				.b4(W2N11D),
				.b5(W2N12D),
				.b6(W2N20D),
				.b7(W2N21D),
				.b8(W2N22D),
				.c(c2D02N)
);

ninexnine_unit ninexnine_unit_6322(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2N00E),
				.b1(W2N01E),
				.b2(W2N02E),
				.b3(W2N10E),
				.b4(W2N11E),
				.b5(W2N12E),
				.b6(W2N20E),
				.b7(W2N21E),
				.b8(W2N22E),
				.c(c2E02N)
);

ninexnine_unit ninexnine_unit_6323(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2N00F),
				.b1(W2N01F),
				.b2(W2N02F),
				.b3(W2N10F),
				.b4(W2N11F),
				.b5(W2N12F),
				.b6(W2N20F),
				.b7(W2N21F),
				.b8(W2N22F),
				.c(c2F02N)
);

assign C202N=c2002N+c2102N+c2202N+c2302N+c2402N+c2502N+c2602N+c2702N+c2802N+c2902N+c2A02N+c2B02N+c2C02N+c2D02N+c2E02N+c2F02N;
assign A202N=(C202N>=0)?1:0;

assign P302N=A202N;

ninexnine_unit ninexnine_unit_6324(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2N000),
				.b1(W2N010),
				.b2(W2N020),
				.b3(W2N100),
				.b4(W2N110),
				.b5(W2N120),
				.b6(W2N200),
				.b7(W2N210),
				.b8(W2N220),
				.c(c2010N)
);

ninexnine_unit ninexnine_unit_6325(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2N001),
				.b1(W2N011),
				.b2(W2N021),
				.b3(W2N101),
				.b4(W2N111),
				.b5(W2N121),
				.b6(W2N201),
				.b7(W2N211),
				.b8(W2N221),
				.c(c2110N)
);

ninexnine_unit ninexnine_unit_6326(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2N002),
				.b1(W2N012),
				.b2(W2N022),
				.b3(W2N102),
				.b4(W2N112),
				.b5(W2N122),
				.b6(W2N202),
				.b7(W2N212),
				.b8(W2N222),
				.c(c2210N)
);

ninexnine_unit ninexnine_unit_6327(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2N003),
				.b1(W2N013),
				.b2(W2N023),
				.b3(W2N103),
				.b4(W2N113),
				.b5(W2N123),
				.b6(W2N203),
				.b7(W2N213),
				.b8(W2N223),
				.c(c2310N)
);

ninexnine_unit ninexnine_unit_6328(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2N004),
				.b1(W2N014),
				.b2(W2N024),
				.b3(W2N104),
				.b4(W2N114),
				.b5(W2N124),
				.b6(W2N204),
				.b7(W2N214),
				.b8(W2N224),
				.c(c2410N)
);

ninexnine_unit ninexnine_unit_6329(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2N005),
				.b1(W2N015),
				.b2(W2N025),
				.b3(W2N105),
				.b4(W2N115),
				.b5(W2N125),
				.b6(W2N205),
				.b7(W2N215),
				.b8(W2N225),
				.c(c2510N)
);

ninexnine_unit ninexnine_unit_6330(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2N006),
				.b1(W2N016),
				.b2(W2N026),
				.b3(W2N106),
				.b4(W2N116),
				.b5(W2N126),
				.b6(W2N206),
				.b7(W2N216),
				.b8(W2N226),
				.c(c2610N)
);

ninexnine_unit ninexnine_unit_6331(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2N007),
				.b1(W2N017),
				.b2(W2N027),
				.b3(W2N107),
				.b4(W2N117),
				.b5(W2N127),
				.b6(W2N207),
				.b7(W2N217),
				.b8(W2N227),
				.c(c2710N)
);

ninexnine_unit ninexnine_unit_6332(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2N008),
				.b1(W2N018),
				.b2(W2N028),
				.b3(W2N108),
				.b4(W2N118),
				.b5(W2N128),
				.b6(W2N208),
				.b7(W2N218),
				.b8(W2N228),
				.c(c2810N)
);

ninexnine_unit ninexnine_unit_6333(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2N009),
				.b1(W2N019),
				.b2(W2N029),
				.b3(W2N109),
				.b4(W2N119),
				.b5(W2N129),
				.b6(W2N209),
				.b7(W2N219),
				.b8(W2N229),
				.c(c2910N)
);

ninexnine_unit ninexnine_unit_6334(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2N00A),
				.b1(W2N01A),
				.b2(W2N02A),
				.b3(W2N10A),
				.b4(W2N11A),
				.b5(W2N12A),
				.b6(W2N20A),
				.b7(W2N21A),
				.b8(W2N22A),
				.c(c2A10N)
);

ninexnine_unit ninexnine_unit_6335(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2N00B),
				.b1(W2N01B),
				.b2(W2N02B),
				.b3(W2N10B),
				.b4(W2N11B),
				.b5(W2N12B),
				.b6(W2N20B),
				.b7(W2N21B),
				.b8(W2N22B),
				.c(c2B10N)
);

ninexnine_unit ninexnine_unit_6336(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2N00C),
				.b1(W2N01C),
				.b2(W2N02C),
				.b3(W2N10C),
				.b4(W2N11C),
				.b5(W2N12C),
				.b6(W2N20C),
				.b7(W2N21C),
				.b8(W2N22C),
				.c(c2C10N)
);

ninexnine_unit ninexnine_unit_6337(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2N00D),
				.b1(W2N01D),
				.b2(W2N02D),
				.b3(W2N10D),
				.b4(W2N11D),
				.b5(W2N12D),
				.b6(W2N20D),
				.b7(W2N21D),
				.b8(W2N22D),
				.c(c2D10N)
);

ninexnine_unit ninexnine_unit_6338(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2N00E),
				.b1(W2N01E),
				.b2(W2N02E),
				.b3(W2N10E),
				.b4(W2N11E),
				.b5(W2N12E),
				.b6(W2N20E),
				.b7(W2N21E),
				.b8(W2N22E),
				.c(c2E10N)
);

ninexnine_unit ninexnine_unit_6339(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2N00F),
				.b1(W2N01F),
				.b2(W2N02F),
				.b3(W2N10F),
				.b4(W2N11F),
				.b5(W2N12F),
				.b6(W2N20F),
				.b7(W2N21F),
				.b8(W2N22F),
				.c(c2F10N)
);

assign C210N=c2010N+c2110N+c2210N+c2310N+c2410N+c2510N+c2610N+c2710N+c2810N+c2910N+c2A10N+c2B10N+c2C10N+c2D10N+c2E10N+c2F10N;
assign A210N=(C210N>=0)?1:0;

assign P310N=A210N;

ninexnine_unit ninexnine_unit_6340(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2N000),
				.b1(W2N010),
				.b2(W2N020),
				.b3(W2N100),
				.b4(W2N110),
				.b5(W2N120),
				.b6(W2N200),
				.b7(W2N210),
				.b8(W2N220),
				.c(c2011N)
);

ninexnine_unit ninexnine_unit_6341(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2N001),
				.b1(W2N011),
				.b2(W2N021),
				.b3(W2N101),
				.b4(W2N111),
				.b5(W2N121),
				.b6(W2N201),
				.b7(W2N211),
				.b8(W2N221),
				.c(c2111N)
);

ninexnine_unit ninexnine_unit_6342(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2N002),
				.b1(W2N012),
				.b2(W2N022),
				.b3(W2N102),
				.b4(W2N112),
				.b5(W2N122),
				.b6(W2N202),
				.b7(W2N212),
				.b8(W2N222),
				.c(c2211N)
);

ninexnine_unit ninexnine_unit_6343(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2N003),
				.b1(W2N013),
				.b2(W2N023),
				.b3(W2N103),
				.b4(W2N113),
				.b5(W2N123),
				.b6(W2N203),
				.b7(W2N213),
				.b8(W2N223),
				.c(c2311N)
);

ninexnine_unit ninexnine_unit_6344(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2N004),
				.b1(W2N014),
				.b2(W2N024),
				.b3(W2N104),
				.b4(W2N114),
				.b5(W2N124),
				.b6(W2N204),
				.b7(W2N214),
				.b8(W2N224),
				.c(c2411N)
);

ninexnine_unit ninexnine_unit_6345(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2N005),
				.b1(W2N015),
				.b2(W2N025),
				.b3(W2N105),
				.b4(W2N115),
				.b5(W2N125),
				.b6(W2N205),
				.b7(W2N215),
				.b8(W2N225),
				.c(c2511N)
);

ninexnine_unit ninexnine_unit_6346(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2N006),
				.b1(W2N016),
				.b2(W2N026),
				.b3(W2N106),
				.b4(W2N116),
				.b5(W2N126),
				.b6(W2N206),
				.b7(W2N216),
				.b8(W2N226),
				.c(c2611N)
);

ninexnine_unit ninexnine_unit_6347(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2N007),
				.b1(W2N017),
				.b2(W2N027),
				.b3(W2N107),
				.b4(W2N117),
				.b5(W2N127),
				.b6(W2N207),
				.b7(W2N217),
				.b8(W2N227),
				.c(c2711N)
);

ninexnine_unit ninexnine_unit_6348(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2N008),
				.b1(W2N018),
				.b2(W2N028),
				.b3(W2N108),
				.b4(W2N118),
				.b5(W2N128),
				.b6(W2N208),
				.b7(W2N218),
				.b8(W2N228),
				.c(c2811N)
);

ninexnine_unit ninexnine_unit_6349(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2N009),
				.b1(W2N019),
				.b2(W2N029),
				.b3(W2N109),
				.b4(W2N119),
				.b5(W2N129),
				.b6(W2N209),
				.b7(W2N219),
				.b8(W2N229),
				.c(c2911N)
);

ninexnine_unit ninexnine_unit_6350(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2N00A),
				.b1(W2N01A),
				.b2(W2N02A),
				.b3(W2N10A),
				.b4(W2N11A),
				.b5(W2N12A),
				.b6(W2N20A),
				.b7(W2N21A),
				.b8(W2N22A),
				.c(c2A11N)
);

ninexnine_unit ninexnine_unit_6351(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2N00B),
				.b1(W2N01B),
				.b2(W2N02B),
				.b3(W2N10B),
				.b4(W2N11B),
				.b5(W2N12B),
				.b6(W2N20B),
				.b7(W2N21B),
				.b8(W2N22B),
				.c(c2B11N)
);

ninexnine_unit ninexnine_unit_6352(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2N00C),
				.b1(W2N01C),
				.b2(W2N02C),
				.b3(W2N10C),
				.b4(W2N11C),
				.b5(W2N12C),
				.b6(W2N20C),
				.b7(W2N21C),
				.b8(W2N22C),
				.c(c2C11N)
);

ninexnine_unit ninexnine_unit_6353(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2N00D),
				.b1(W2N01D),
				.b2(W2N02D),
				.b3(W2N10D),
				.b4(W2N11D),
				.b5(W2N12D),
				.b6(W2N20D),
				.b7(W2N21D),
				.b8(W2N22D),
				.c(c2D11N)
);

ninexnine_unit ninexnine_unit_6354(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2N00E),
				.b1(W2N01E),
				.b2(W2N02E),
				.b3(W2N10E),
				.b4(W2N11E),
				.b5(W2N12E),
				.b6(W2N20E),
				.b7(W2N21E),
				.b8(W2N22E),
				.c(c2E11N)
);

ninexnine_unit ninexnine_unit_6355(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2N00F),
				.b1(W2N01F),
				.b2(W2N02F),
				.b3(W2N10F),
				.b4(W2N11F),
				.b5(W2N12F),
				.b6(W2N20F),
				.b7(W2N21F),
				.b8(W2N22F),
				.c(c2F11N)
);

assign C211N=c2011N+c2111N+c2211N+c2311N+c2411N+c2511N+c2611N+c2711N+c2811N+c2911N+c2A11N+c2B11N+c2C11N+c2D11N+c2E11N+c2F11N;
assign A211N=(C211N>=0)?1:0;

assign P311N=A211N;

ninexnine_unit ninexnine_unit_6356(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2N000),
				.b1(W2N010),
				.b2(W2N020),
				.b3(W2N100),
				.b4(W2N110),
				.b5(W2N120),
				.b6(W2N200),
				.b7(W2N210),
				.b8(W2N220),
				.c(c2012N)
);

ninexnine_unit ninexnine_unit_6357(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2N001),
				.b1(W2N011),
				.b2(W2N021),
				.b3(W2N101),
				.b4(W2N111),
				.b5(W2N121),
				.b6(W2N201),
				.b7(W2N211),
				.b8(W2N221),
				.c(c2112N)
);

ninexnine_unit ninexnine_unit_6358(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2N002),
				.b1(W2N012),
				.b2(W2N022),
				.b3(W2N102),
				.b4(W2N112),
				.b5(W2N122),
				.b6(W2N202),
				.b7(W2N212),
				.b8(W2N222),
				.c(c2212N)
);

ninexnine_unit ninexnine_unit_6359(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2N003),
				.b1(W2N013),
				.b2(W2N023),
				.b3(W2N103),
				.b4(W2N113),
				.b5(W2N123),
				.b6(W2N203),
				.b7(W2N213),
				.b8(W2N223),
				.c(c2312N)
);

ninexnine_unit ninexnine_unit_6360(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2N004),
				.b1(W2N014),
				.b2(W2N024),
				.b3(W2N104),
				.b4(W2N114),
				.b5(W2N124),
				.b6(W2N204),
				.b7(W2N214),
				.b8(W2N224),
				.c(c2412N)
);

ninexnine_unit ninexnine_unit_6361(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2N005),
				.b1(W2N015),
				.b2(W2N025),
				.b3(W2N105),
				.b4(W2N115),
				.b5(W2N125),
				.b6(W2N205),
				.b7(W2N215),
				.b8(W2N225),
				.c(c2512N)
);

ninexnine_unit ninexnine_unit_6362(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2N006),
				.b1(W2N016),
				.b2(W2N026),
				.b3(W2N106),
				.b4(W2N116),
				.b5(W2N126),
				.b6(W2N206),
				.b7(W2N216),
				.b8(W2N226),
				.c(c2612N)
);

ninexnine_unit ninexnine_unit_6363(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2N007),
				.b1(W2N017),
				.b2(W2N027),
				.b3(W2N107),
				.b4(W2N117),
				.b5(W2N127),
				.b6(W2N207),
				.b7(W2N217),
				.b8(W2N227),
				.c(c2712N)
);

ninexnine_unit ninexnine_unit_6364(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2N008),
				.b1(W2N018),
				.b2(W2N028),
				.b3(W2N108),
				.b4(W2N118),
				.b5(W2N128),
				.b6(W2N208),
				.b7(W2N218),
				.b8(W2N228),
				.c(c2812N)
);

ninexnine_unit ninexnine_unit_6365(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2N009),
				.b1(W2N019),
				.b2(W2N029),
				.b3(W2N109),
				.b4(W2N119),
				.b5(W2N129),
				.b6(W2N209),
				.b7(W2N219),
				.b8(W2N229),
				.c(c2912N)
);

ninexnine_unit ninexnine_unit_6366(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2N00A),
				.b1(W2N01A),
				.b2(W2N02A),
				.b3(W2N10A),
				.b4(W2N11A),
				.b5(W2N12A),
				.b6(W2N20A),
				.b7(W2N21A),
				.b8(W2N22A),
				.c(c2A12N)
);

ninexnine_unit ninexnine_unit_6367(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2N00B),
				.b1(W2N01B),
				.b2(W2N02B),
				.b3(W2N10B),
				.b4(W2N11B),
				.b5(W2N12B),
				.b6(W2N20B),
				.b7(W2N21B),
				.b8(W2N22B),
				.c(c2B12N)
);

ninexnine_unit ninexnine_unit_6368(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2N00C),
				.b1(W2N01C),
				.b2(W2N02C),
				.b3(W2N10C),
				.b4(W2N11C),
				.b5(W2N12C),
				.b6(W2N20C),
				.b7(W2N21C),
				.b8(W2N22C),
				.c(c2C12N)
);

ninexnine_unit ninexnine_unit_6369(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2N00D),
				.b1(W2N01D),
				.b2(W2N02D),
				.b3(W2N10D),
				.b4(W2N11D),
				.b5(W2N12D),
				.b6(W2N20D),
				.b7(W2N21D),
				.b8(W2N22D),
				.c(c2D12N)
);

ninexnine_unit ninexnine_unit_6370(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2N00E),
				.b1(W2N01E),
				.b2(W2N02E),
				.b3(W2N10E),
				.b4(W2N11E),
				.b5(W2N12E),
				.b6(W2N20E),
				.b7(W2N21E),
				.b8(W2N22E),
				.c(c2E12N)
);

ninexnine_unit ninexnine_unit_6371(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2N00F),
				.b1(W2N01F),
				.b2(W2N02F),
				.b3(W2N10F),
				.b4(W2N11F),
				.b5(W2N12F),
				.b6(W2N20F),
				.b7(W2N21F),
				.b8(W2N22F),
				.c(c2F12N)
);

assign C212N=c2012N+c2112N+c2212N+c2312N+c2412N+c2512N+c2612N+c2712N+c2812N+c2912N+c2A12N+c2B12N+c2C12N+c2D12N+c2E12N+c2F12N;
assign A212N=(C212N>=0)?1:0;

assign P312N=A212N;

ninexnine_unit ninexnine_unit_6372(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2N000),
				.b1(W2N010),
				.b2(W2N020),
				.b3(W2N100),
				.b4(W2N110),
				.b5(W2N120),
				.b6(W2N200),
				.b7(W2N210),
				.b8(W2N220),
				.c(c2020N)
);

ninexnine_unit ninexnine_unit_6373(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2N001),
				.b1(W2N011),
				.b2(W2N021),
				.b3(W2N101),
				.b4(W2N111),
				.b5(W2N121),
				.b6(W2N201),
				.b7(W2N211),
				.b8(W2N221),
				.c(c2120N)
);

ninexnine_unit ninexnine_unit_6374(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2N002),
				.b1(W2N012),
				.b2(W2N022),
				.b3(W2N102),
				.b4(W2N112),
				.b5(W2N122),
				.b6(W2N202),
				.b7(W2N212),
				.b8(W2N222),
				.c(c2220N)
);

ninexnine_unit ninexnine_unit_6375(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2N003),
				.b1(W2N013),
				.b2(W2N023),
				.b3(W2N103),
				.b4(W2N113),
				.b5(W2N123),
				.b6(W2N203),
				.b7(W2N213),
				.b8(W2N223),
				.c(c2320N)
);

ninexnine_unit ninexnine_unit_6376(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2N004),
				.b1(W2N014),
				.b2(W2N024),
				.b3(W2N104),
				.b4(W2N114),
				.b5(W2N124),
				.b6(W2N204),
				.b7(W2N214),
				.b8(W2N224),
				.c(c2420N)
);

ninexnine_unit ninexnine_unit_6377(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2N005),
				.b1(W2N015),
				.b2(W2N025),
				.b3(W2N105),
				.b4(W2N115),
				.b5(W2N125),
				.b6(W2N205),
				.b7(W2N215),
				.b8(W2N225),
				.c(c2520N)
);

ninexnine_unit ninexnine_unit_6378(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2N006),
				.b1(W2N016),
				.b2(W2N026),
				.b3(W2N106),
				.b4(W2N116),
				.b5(W2N126),
				.b6(W2N206),
				.b7(W2N216),
				.b8(W2N226),
				.c(c2620N)
);

ninexnine_unit ninexnine_unit_6379(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2N007),
				.b1(W2N017),
				.b2(W2N027),
				.b3(W2N107),
				.b4(W2N117),
				.b5(W2N127),
				.b6(W2N207),
				.b7(W2N217),
				.b8(W2N227),
				.c(c2720N)
);

ninexnine_unit ninexnine_unit_6380(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2N008),
				.b1(W2N018),
				.b2(W2N028),
				.b3(W2N108),
				.b4(W2N118),
				.b5(W2N128),
				.b6(W2N208),
				.b7(W2N218),
				.b8(W2N228),
				.c(c2820N)
);

ninexnine_unit ninexnine_unit_6381(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2N009),
				.b1(W2N019),
				.b2(W2N029),
				.b3(W2N109),
				.b4(W2N119),
				.b5(W2N129),
				.b6(W2N209),
				.b7(W2N219),
				.b8(W2N229),
				.c(c2920N)
);

ninexnine_unit ninexnine_unit_6382(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2N00A),
				.b1(W2N01A),
				.b2(W2N02A),
				.b3(W2N10A),
				.b4(W2N11A),
				.b5(W2N12A),
				.b6(W2N20A),
				.b7(W2N21A),
				.b8(W2N22A),
				.c(c2A20N)
);

ninexnine_unit ninexnine_unit_6383(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2N00B),
				.b1(W2N01B),
				.b2(W2N02B),
				.b3(W2N10B),
				.b4(W2N11B),
				.b5(W2N12B),
				.b6(W2N20B),
				.b7(W2N21B),
				.b8(W2N22B),
				.c(c2B20N)
);

ninexnine_unit ninexnine_unit_6384(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2N00C),
				.b1(W2N01C),
				.b2(W2N02C),
				.b3(W2N10C),
				.b4(W2N11C),
				.b5(W2N12C),
				.b6(W2N20C),
				.b7(W2N21C),
				.b8(W2N22C),
				.c(c2C20N)
);

ninexnine_unit ninexnine_unit_6385(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2N00D),
				.b1(W2N01D),
				.b2(W2N02D),
				.b3(W2N10D),
				.b4(W2N11D),
				.b5(W2N12D),
				.b6(W2N20D),
				.b7(W2N21D),
				.b8(W2N22D),
				.c(c2D20N)
);

ninexnine_unit ninexnine_unit_6386(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2N00E),
				.b1(W2N01E),
				.b2(W2N02E),
				.b3(W2N10E),
				.b4(W2N11E),
				.b5(W2N12E),
				.b6(W2N20E),
				.b7(W2N21E),
				.b8(W2N22E),
				.c(c2E20N)
);

ninexnine_unit ninexnine_unit_6387(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2N00F),
				.b1(W2N01F),
				.b2(W2N02F),
				.b3(W2N10F),
				.b4(W2N11F),
				.b5(W2N12F),
				.b6(W2N20F),
				.b7(W2N21F),
				.b8(W2N22F),
				.c(c2F20N)
);

assign C220N=c2020N+c2120N+c2220N+c2320N+c2420N+c2520N+c2620N+c2720N+c2820N+c2920N+c2A20N+c2B20N+c2C20N+c2D20N+c2E20N+c2F20N;
assign A220N=(C220N>=0)?1:0;

assign P320N=A220N;

ninexnine_unit ninexnine_unit_6388(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2N000),
				.b1(W2N010),
				.b2(W2N020),
				.b3(W2N100),
				.b4(W2N110),
				.b5(W2N120),
				.b6(W2N200),
				.b7(W2N210),
				.b8(W2N220),
				.c(c2021N)
);

ninexnine_unit ninexnine_unit_6389(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2N001),
				.b1(W2N011),
				.b2(W2N021),
				.b3(W2N101),
				.b4(W2N111),
				.b5(W2N121),
				.b6(W2N201),
				.b7(W2N211),
				.b8(W2N221),
				.c(c2121N)
);

ninexnine_unit ninexnine_unit_6390(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2N002),
				.b1(W2N012),
				.b2(W2N022),
				.b3(W2N102),
				.b4(W2N112),
				.b5(W2N122),
				.b6(W2N202),
				.b7(W2N212),
				.b8(W2N222),
				.c(c2221N)
);

ninexnine_unit ninexnine_unit_6391(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2N003),
				.b1(W2N013),
				.b2(W2N023),
				.b3(W2N103),
				.b4(W2N113),
				.b5(W2N123),
				.b6(W2N203),
				.b7(W2N213),
				.b8(W2N223),
				.c(c2321N)
);

ninexnine_unit ninexnine_unit_6392(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2N004),
				.b1(W2N014),
				.b2(W2N024),
				.b3(W2N104),
				.b4(W2N114),
				.b5(W2N124),
				.b6(W2N204),
				.b7(W2N214),
				.b8(W2N224),
				.c(c2421N)
);

ninexnine_unit ninexnine_unit_6393(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2N005),
				.b1(W2N015),
				.b2(W2N025),
				.b3(W2N105),
				.b4(W2N115),
				.b5(W2N125),
				.b6(W2N205),
				.b7(W2N215),
				.b8(W2N225),
				.c(c2521N)
);

ninexnine_unit ninexnine_unit_6394(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2N006),
				.b1(W2N016),
				.b2(W2N026),
				.b3(W2N106),
				.b4(W2N116),
				.b5(W2N126),
				.b6(W2N206),
				.b7(W2N216),
				.b8(W2N226),
				.c(c2621N)
);

ninexnine_unit ninexnine_unit_6395(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2N007),
				.b1(W2N017),
				.b2(W2N027),
				.b3(W2N107),
				.b4(W2N117),
				.b5(W2N127),
				.b6(W2N207),
				.b7(W2N217),
				.b8(W2N227),
				.c(c2721N)
);

ninexnine_unit ninexnine_unit_6396(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2N008),
				.b1(W2N018),
				.b2(W2N028),
				.b3(W2N108),
				.b4(W2N118),
				.b5(W2N128),
				.b6(W2N208),
				.b7(W2N218),
				.b8(W2N228),
				.c(c2821N)
);

ninexnine_unit ninexnine_unit_6397(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2N009),
				.b1(W2N019),
				.b2(W2N029),
				.b3(W2N109),
				.b4(W2N119),
				.b5(W2N129),
				.b6(W2N209),
				.b7(W2N219),
				.b8(W2N229),
				.c(c2921N)
);

ninexnine_unit ninexnine_unit_6398(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2N00A),
				.b1(W2N01A),
				.b2(W2N02A),
				.b3(W2N10A),
				.b4(W2N11A),
				.b5(W2N12A),
				.b6(W2N20A),
				.b7(W2N21A),
				.b8(W2N22A),
				.c(c2A21N)
);

ninexnine_unit ninexnine_unit_6399(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2N00B),
				.b1(W2N01B),
				.b2(W2N02B),
				.b3(W2N10B),
				.b4(W2N11B),
				.b5(W2N12B),
				.b6(W2N20B),
				.b7(W2N21B),
				.b8(W2N22B),
				.c(c2B21N)
);

ninexnine_unit ninexnine_unit_6400(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2N00C),
				.b1(W2N01C),
				.b2(W2N02C),
				.b3(W2N10C),
				.b4(W2N11C),
				.b5(W2N12C),
				.b6(W2N20C),
				.b7(W2N21C),
				.b8(W2N22C),
				.c(c2C21N)
);

ninexnine_unit ninexnine_unit_6401(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2N00D),
				.b1(W2N01D),
				.b2(W2N02D),
				.b3(W2N10D),
				.b4(W2N11D),
				.b5(W2N12D),
				.b6(W2N20D),
				.b7(W2N21D),
				.b8(W2N22D),
				.c(c2D21N)
);

ninexnine_unit ninexnine_unit_6402(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2N00E),
				.b1(W2N01E),
				.b2(W2N02E),
				.b3(W2N10E),
				.b4(W2N11E),
				.b5(W2N12E),
				.b6(W2N20E),
				.b7(W2N21E),
				.b8(W2N22E),
				.c(c2E21N)
);

ninexnine_unit ninexnine_unit_6403(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2N00F),
				.b1(W2N01F),
				.b2(W2N02F),
				.b3(W2N10F),
				.b4(W2N11F),
				.b5(W2N12F),
				.b6(W2N20F),
				.b7(W2N21F),
				.b8(W2N22F),
				.c(c2F21N)
);

assign C221N=c2021N+c2121N+c2221N+c2321N+c2421N+c2521N+c2621N+c2721N+c2821N+c2921N+c2A21N+c2B21N+c2C21N+c2D21N+c2E21N+c2F21N;
assign A221N=(C221N>=0)?1:0;

assign P321N=A221N;

ninexnine_unit ninexnine_unit_6404(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2N000),
				.b1(W2N010),
				.b2(W2N020),
				.b3(W2N100),
				.b4(W2N110),
				.b5(W2N120),
				.b6(W2N200),
				.b7(W2N210),
				.b8(W2N220),
				.c(c2022N)
);

ninexnine_unit ninexnine_unit_6405(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2N001),
				.b1(W2N011),
				.b2(W2N021),
				.b3(W2N101),
				.b4(W2N111),
				.b5(W2N121),
				.b6(W2N201),
				.b7(W2N211),
				.b8(W2N221),
				.c(c2122N)
);

ninexnine_unit ninexnine_unit_6406(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2N002),
				.b1(W2N012),
				.b2(W2N022),
				.b3(W2N102),
				.b4(W2N112),
				.b5(W2N122),
				.b6(W2N202),
				.b7(W2N212),
				.b8(W2N222),
				.c(c2222N)
);

ninexnine_unit ninexnine_unit_6407(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2N003),
				.b1(W2N013),
				.b2(W2N023),
				.b3(W2N103),
				.b4(W2N113),
				.b5(W2N123),
				.b6(W2N203),
				.b7(W2N213),
				.b8(W2N223),
				.c(c2322N)
);

ninexnine_unit ninexnine_unit_6408(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2N004),
				.b1(W2N014),
				.b2(W2N024),
				.b3(W2N104),
				.b4(W2N114),
				.b5(W2N124),
				.b6(W2N204),
				.b7(W2N214),
				.b8(W2N224),
				.c(c2422N)
);

ninexnine_unit ninexnine_unit_6409(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2N005),
				.b1(W2N015),
				.b2(W2N025),
				.b3(W2N105),
				.b4(W2N115),
				.b5(W2N125),
				.b6(W2N205),
				.b7(W2N215),
				.b8(W2N225),
				.c(c2522N)
);

ninexnine_unit ninexnine_unit_6410(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2N006),
				.b1(W2N016),
				.b2(W2N026),
				.b3(W2N106),
				.b4(W2N116),
				.b5(W2N126),
				.b6(W2N206),
				.b7(W2N216),
				.b8(W2N226),
				.c(c2622N)
);

ninexnine_unit ninexnine_unit_6411(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2N007),
				.b1(W2N017),
				.b2(W2N027),
				.b3(W2N107),
				.b4(W2N117),
				.b5(W2N127),
				.b6(W2N207),
				.b7(W2N217),
				.b8(W2N227),
				.c(c2722N)
);

ninexnine_unit ninexnine_unit_6412(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2N008),
				.b1(W2N018),
				.b2(W2N028),
				.b3(W2N108),
				.b4(W2N118),
				.b5(W2N128),
				.b6(W2N208),
				.b7(W2N218),
				.b8(W2N228),
				.c(c2822N)
);

ninexnine_unit ninexnine_unit_6413(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2N009),
				.b1(W2N019),
				.b2(W2N029),
				.b3(W2N109),
				.b4(W2N119),
				.b5(W2N129),
				.b6(W2N209),
				.b7(W2N219),
				.b8(W2N229),
				.c(c2922N)
);

ninexnine_unit ninexnine_unit_6414(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2N00A),
				.b1(W2N01A),
				.b2(W2N02A),
				.b3(W2N10A),
				.b4(W2N11A),
				.b5(W2N12A),
				.b6(W2N20A),
				.b7(W2N21A),
				.b8(W2N22A),
				.c(c2A22N)
);

ninexnine_unit ninexnine_unit_6415(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2N00B),
				.b1(W2N01B),
				.b2(W2N02B),
				.b3(W2N10B),
				.b4(W2N11B),
				.b5(W2N12B),
				.b6(W2N20B),
				.b7(W2N21B),
				.b8(W2N22B),
				.c(c2B22N)
);

ninexnine_unit ninexnine_unit_6416(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2N00C),
				.b1(W2N01C),
				.b2(W2N02C),
				.b3(W2N10C),
				.b4(W2N11C),
				.b5(W2N12C),
				.b6(W2N20C),
				.b7(W2N21C),
				.b8(W2N22C),
				.c(c2C22N)
);

ninexnine_unit ninexnine_unit_6417(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2N00D),
				.b1(W2N01D),
				.b2(W2N02D),
				.b3(W2N10D),
				.b4(W2N11D),
				.b5(W2N12D),
				.b6(W2N20D),
				.b7(W2N21D),
				.b8(W2N22D),
				.c(c2D22N)
);

ninexnine_unit ninexnine_unit_6418(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2N00E),
				.b1(W2N01E),
				.b2(W2N02E),
				.b3(W2N10E),
				.b4(W2N11E),
				.b5(W2N12E),
				.b6(W2N20E),
				.b7(W2N21E),
				.b8(W2N22E),
				.c(c2E22N)
);

ninexnine_unit ninexnine_unit_6419(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2N00F),
				.b1(W2N01F),
				.b2(W2N02F),
				.b3(W2N10F),
				.b4(W2N11F),
				.b5(W2N12F),
				.b6(W2N20F),
				.b7(W2N21F),
				.b8(W2N22F),
				.c(c2F22N)
);

assign C222N=c2022N+c2122N+c2222N+c2322N+c2422N+c2522N+c2622N+c2722N+c2822N+c2922N+c2A22N+c2B22N+c2C22N+c2D22N+c2E22N+c2F22N;
assign A222N=(C222N>=0)?1:0;

assign P322N=A222N;

ninexnine_unit ninexnine_unit_6420(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2O000),
				.b1(W2O010),
				.b2(W2O020),
				.b3(W2O100),
				.b4(W2O110),
				.b5(W2O120),
				.b6(W2O200),
				.b7(W2O210),
				.b8(W2O220),
				.c(c2000O)
);

ninexnine_unit ninexnine_unit_6421(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2O001),
				.b1(W2O011),
				.b2(W2O021),
				.b3(W2O101),
				.b4(W2O111),
				.b5(W2O121),
				.b6(W2O201),
				.b7(W2O211),
				.b8(W2O221),
				.c(c2100O)
);

ninexnine_unit ninexnine_unit_6422(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2O002),
				.b1(W2O012),
				.b2(W2O022),
				.b3(W2O102),
				.b4(W2O112),
				.b5(W2O122),
				.b6(W2O202),
				.b7(W2O212),
				.b8(W2O222),
				.c(c2200O)
);

ninexnine_unit ninexnine_unit_6423(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2O003),
				.b1(W2O013),
				.b2(W2O023),
				.b3(W2O103),
				.b4(W2O113),
				.b5(W2O123),
				.b6(W2O203),
				.b7(W2O213),
				.b8(W2O223),
				.c(c2300O)
);

ninexnine_unit ninexnine_unit_6424(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2O004),
				.b1(W2O014),
				.b2(W2O024),
				.b3(W2O104),
				.b4(W2O114),
				.b5(W2O124),
				.b6(W2O204),
				.b7(W2O214),
				.b8(W2O224),
				.c(c2400O)
);

ninexnine_unit ninexnine_unit_6425(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2O005),
				.b1(W2O015),
				.b2(W2O025),
				.b3(W2O105),
				.b4(W2O115),
				.b5(W2O125),
				.b6(W2O205),
				.b7(W2O215),
				.b8(W2O225),
				.c(c2500O)
);

ninexnine_unit ninexnine_unit_6426(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2O006),
				.b1(W2O016),
				.b2(W2O026),
				.b3(W2O106),
				.b4(W2O116),
				.b5(W2O126),
				.b6(W2O206),
				.b7(W2O216),
				.b8(W2O226),
				.c(c2600O)
);

ninexnine_unit ninexnine_unit_6427(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2O007),
				.b1(W2O017),
				.b2(W2O027),
				.b3(W2O107),
				.b4(W2O117),
				.b5(W2O127),
				.b6(W2O207),
				.b7(W2O217),
				.b8(W2O227),
				.c(c2700O)
);

ninexnine_unit ninexnine_unit_6428(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2O008),
				.b1(W2O018),
				.b2(W2O028),
				.b3(W2O108),
				.b4(W2O118),
				.b5(W2O128),
				.b6(W2O208),
				.b7(W2O218),
				.b8(W2O228),
				.c(c2800O)
);

ninexnine_unit ninexnine_unit_6429(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2O009),
				.b1(W2O019),
				.b2(W2O029),
				.b3(W2O109),
				.b4(W2O119),
				.b5(W2O129),
				.b6(W2O209),
				.b7(W2O219),
				.b8(W2O229),
				.c(c2900O)
);

ninexnine_unit ninexnine_unit_6430(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2O00A),
				.b1(W2O01A),
				.b2(W2O02A),
				.b3(W2O10A),
				.b4(W2O11A),
				.b5(W2O12A),
				.b6(W2O20A),
				.b7(W2O21A),
				.b8(W2O22A),
				.c(c2A00O)
);

ninexnine_unit ninexnine_unit_6431(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2O00B),
				.b1(W2O01B),
				.b2(W2O02B),
				.b3(W2O10B),
				.b4(W2O11B),
				.b5(W2O12B),
				.b6(W2O20B),
				.b7(W2O21B),
				.b8(W2O22B),
				.c(c2B00O)
);

ninexnine_unit ninexnine_unit_6432(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2O00C),
				.b1(W2O01C),
				.b2(W2O02C),
				.b3(W2O10C),
				.b4(W2O11C),
				.b5(W2O12C),
				.b6(W2O20C),
				.b7(W2O21C),
				.b8(W2O22C),
				.c(c2C00O)
);

ninexnine_unit ninexnine_unit_6433(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2O00D),
				.b1(W2O01D),
				.b2(W2O02D),
				.b3(W2O10D),
				.b4(W2O11D),
				.b5(W2O12D),
				.b6(W2O20D),
				.b7(W2O21D),
				.b8(W2O22D),
				.c(c2D00O)
);

ninexnine_unit ninexnine_unit_6434(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2O00E),
				.b1(W2O01E),
				.b2(W2O02E),
				.b3(W2O10E),
				.b4(W2O11E),
				.b5(W2O12E),
				.b6(W2O20E),
				.b7(W2O21E),
				.b8(W2O22E),
				.c(c2E00O)
);

ninexnine_unit ninexnine_unit_6435(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2O00F),
				.b1(W2O01F),
				.b2(W2O02F),
				.b3(W2O10F),
				.b4(W2O11F),
				.b5(W2O12F),
				.b6(W2O20F),
				.b7(W2O21F),
				.b8(W2O22F),
				.c(c2F00O)
);

assign C200O=c2000O+c2100O+c2200O+c2300O+c2400O+c2500O+c2600O+c2700O+c2800O+c2900O+c2A00O+c2B00O+c2C00O+c2D00O+c2E00O+c2F00O;
assign A200O=(C200O>=0)?1:0;

assign P300O=A200O;

ninexnine_unit ninexnine_unit_6436(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2O000),
				.b1(W2O010),
				.b2(W2O020),
				.b3(W2O100),
				.b4(W2O110),
				.b5(W2O120),
				.b6(W2O200),
				.b7(W2O210),
				.b8(W2O220),
				.c(c2001O)
);

ninexnine_unit ninexnine_unit_6437(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2O001),
				.b1(W2O011),
				.b2(W2O021),
				.b3(W2O101),
				.b4(W2O111),
				.b5(W2O121),
				.b6(W2O201),
				.b7(W2O211),
				.b8(W2O221),
				.c(c2101O)
);

ninexnine_unit ninexnine_unit_6438(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2O002),
				.b1(W2O012),
				.b2(W2O022),
				.b3(W2O102),
				.b4(W2O112),
				.b5(W2O122),
				.b6(W2O202),
				.b7(W2O212),
				.b8(W2O222),
				.c(c2201O)
);

ninexnine_unit ninexnine_unit_6439(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2O003),
				.b1(W2O013),
				.b2(W2O023),
				.b3(W2O103),
				.b4(W2O113),
				.b5(W2O123),
				.b6(W2O203),
				.b7(W2O213),
				.b8(W2O223),
				.c(c2301O)
);

ninexnine_unit ninexnine_unit_6440(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2O004),
				.b1(W2O014),
				.b2(W2O024),
				.b3(W2O104),
				.b4(W2O114),
				.b5(W2O124),
				.b6(W2O204),
				.b7(W2O214),
				.b8(W2O224),
				.c(c2401O)
);

ninexnine_unit ninexnine_unit_6441(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2O005),
				.b1(W2O015),
				.b2(W2O025),
				.b3(W2O105),
				.b4(W2O115),
				.b5(W2O125),
				.b6(W2O205),
				.b7(W2O215),
				.b8(W2O225),
				.c(c2501O)
);

ninexnine_unit ninexnine_unit_6442(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2O006),
				.b1(W2O016),
				.b2(W2O026),
				.b3(W2O106),
				.b4(W2O116),
				.b5(W2O126),
				.b6(W2O206),
				.b7(W2O216),
				.b8(W2O226),
				.c(c2601O)
);

ninexnine_unit ninexnine_unit_6443(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2O007),
				.b1(W2O017),
				.b2(W2O027),
				.b3(W2O107),
				.b4(W2O117),
				.b5(W2O127),
				.b6(W2O207),
				.b7(W2O217),
				.b8(W2O227),
				.c(c2701O)
);

ninexnine_unit ninexnine_unit_6444(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2O008),
				.b1(W2O018),
				.b2(W2O028),
				.b3(W2O108),
				.b4(W2O118),
				.b5(W2O128),
				.b6(W2O208),
				.b7(W2O218),
				.b8(W2O228),
				.c(c2801O)
);

ninexnine_unit ninexnine_unit_6445(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2O009),
				.b1(W2O019),
				.b2(W2O029),
				.b3(W2O109),
				.b4(W2O119),
				.b5(W2O129),
				.b6(W2O209),
				.b7(W2O219),
				.b8(W2O229),
				.c(c2901O)
);

ninexnine_unit ninexnine_unit_6446(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2O00A),
				.b1(W2O01A),
				.b2(W2O02A),
				.b3(W2O10A),
				.b4(W2O11A),
				.b5(W2O12A),
				.b6(W2O20A),
				.b7(W2O21A),
				.b8(W2O22A),
				.c(c2A01O)
);

ninexnine_unit ninexnine_unit_6447(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2O00B),
				.b1(W2O01B),
				.b2(W2O02B),
				.b3(W2O10B),
				.b4(W2O11B),
				.b5(W2O12B),
				.b6(W2O20B),
				.b7(W2O21B),
				.b8(W2O22B),
				.c(c2B01O)
);

ninexnine_unit ninexnine_unit_6448(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2O00C),
				.b1(W2O01C),
				.b2(W2O02C),
				.b3(W2O10C),
				.b4(W2O11C),
				.b5(W2O12C),
				.b6(W2O20C),
				.b7(W2O21C),
				.b8(W2O22C),
				.c(c2C01O)
);

ninexnine_unit ninexnine_unit_6449(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2O00D),
				.b1(W2O01D),
				.b2(W2O02D),
				.b3(W2O10D),
				.b4(W2O11D),
				.b5(W2O12D),
				.b6(W2O20D),
				.b7(W2O21D),
				.b8(W2O22D),
				.c(c2D01O)
);

ninexnine_unit ninexnine_unit_6450(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2O00E),
				.b1(W2O01E),
				.b2(W2O02E),
				.b3(W2O10E),
				.b4(W2O11E),
				.b5(W2O12E),
				.b6(W2O20E),
				.b7(W2O21E),
				.b8(W2O22E),
				.c(c2E01O)
);

ninexnine_unit ninexnine_unit_6451(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2O00F),
				.b1(W2O01F),
				.b2(W2O02F),
				.b3(W2O10F),
				.b4(W2O11F),
				.b5(W2O12F),
				.b6(W2O20F),
				.b7(W2O21F),
				.b8(W2O22F),
				.c(c2F01O)
);

assign C201O=c2001O+c2101O+c2201O+c2301O+c2401O+c2501O+c2601O+c2701O+c2801O+c2901O+c2A01O+c2B01O+c2C01O+c2D01O+c2E01O+c2F01O;
assign A201O=(C201O>=0)?1:0;

assign P301O=A201O;

ninexnine_unit ninexnine_unit_6452(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2O000),
				.b1(W2O010),
				.b2(W2O020),
				.b3(W2O100),
				.b4(W2O110),
				.b5(W2O120),
				.b6(W2O200),
				.b7(W2O210),
				.b8(W2O220),
				.c(c2002O)
);

ninexnine_unit ninexnine_unit_6453(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2O001),
				.b1(W2O011),
				.b2(W2O021),
				.b3(W2O101),
				.b4(W2O111),
				.b5(W2O121),
				.b6(W2O201),
				.b7(W2O211),
				.b8(W2O221),
				.c(c2102O)
);

ninexnine_unit ninexnine_unit_6454(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2O002),
				.b1(W2O012),
				.b2(W2O022),
				.b3(W2O102),
				.b4(W2O112),
				.b5(W2O122),
				.b6(W2O202),
				.b7(W2O212),
				.b8(W2O222),
				.c(c2202O)
);

ninexnine_unit ninexnine_unit_6455(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2O003),
				.b1(W2O013),
				.b2(W2O023),
				.b3(W2O103),
				.b4(W2O113),
				.b5(W2O123),
				.b6(W2O203),
				.b7(W2O213),
				.b8(W2O223),
				.c(c2302O)
);

ninexnine_unit ninexnine_unit_6456(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2O004),
				.b1(W2O014),
				.b2(W2O024),
				.b3(W2O104),
				.b4(W2O114),
				.b5(W2O124),
				.b6(W2O204),
				.b7(W2O214),
				.b8(W2O224),
				.c(c2402O)
);

ninexnine_unit ninexnine_unit_6457(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2O005),
				.b1(W2O015),
				.b2(W2O025),
				.b3(W2O105),
				.b4(W2O115),
				.b5(W2O125),
				.b6(W2O205),
				.b7(W2O215),
				.b8(W2O225),
				.c(c2502O)
);

ninexnine_unit ninexnine_unit_6458(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2O006),
				.b1(W2O016),
				.b2(W2O026),
				.b3(W2O106),
				.b4(W2O116),
				.b5(W2O126),
				.b6(W2O206),
				.b7(W2O216),
				.b8(W2O226),
				.c(c2602O)
);

ninexnine_unit ninexnine_unit_6459(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2O007),
				.b1(W2O017),
				.b2(W2O027),
				.b3(W2O107),
				.b4(W2O117),
				.b5(W2O127),
				.b6(W2O207),
				.b7(W2O217),
				.b8(W2O227),
				.c(c2702O)
);

ninexnine_unit ninexnine_unit_6460(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2O008),
				.b1(W2O018),
				.b2(W2O028),
				.b3(W2O108),
				.b4(W2O118),
				.b5(W2O128),
				.b6(W2O208),
				.b7(W2O218),
				.b8(W2O228),
				.c(c2802O)
);

ninexnine_unit ninexnine_unit_6461(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2O009),
				.b1(W2O019),
				.b2(W2O029),
				.b3(W2O109),
				.b4(W2O119),
				.b5(W2O129),
				.b6(W2O209),
				.b7(W2O219),
				.b8(W2O229),
				.c(c2902O)
);

ninexnine_unit ninexnine_unit_6462(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2O00A),
				.b1(W2O01A),
				.b2(W2O02A),
				.b3(W2O10A),
				.b4(W2O11A),
				.b5(W2O12A),
				.b6(W2O20A),
				.b7(W2O21A),
				.b8(W2O22A),
				.c(c2A02O)
);

ninexnine_unit ninexnine_unit_6463(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2O00B),
				.b1(W2O01B),
				.b2(W2O02B),
				.b3(W2O10B),
				.b4(W2O11B),
				.b5(W2O12B),
				.b6(W2O20B),
				.b7(W2O21B),
				.b8(W2O22B),
				.c(c2B02O)
);

ninexnine_unit ninexnine_unit_6464(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2O00C),
				.b1(W2O01C),
				.b2(W2O02C),
				.b3(W2O10C),
				.b4(W2O11C),
				.b5(W2O12C),
				.b6(W2O20C),
				.b7(W2O21C),
				.b8(W2O22C),
				.c(c2C02O)
);

ninexnine_unit ninexnine_unit_6465(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2O00D),
				.b1(W2O01D),
				.b2(W2O02D),
				.b3(W2O10D),
				.b4(W2O11D),
				.b5(W2O12D),
				.b6(W2O20D),
				.b7(W2O21D),
				.b8(W2O22D),
				.c(c2D02O)
);

ninexnine_unit ninexnine_unit_6466(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2O00E),
				.b1(W2O01E),
				.b2(W2O02E),
				.b3(W2O10E),
				.b4(W2O11E),
				.b5(W2O12E),
				.b6(W2O20E),
				.b7(W2O21E),
				.b8(W2O22E),
				.c(c2E02O)
);

ninexnine_unit ninexnine_unit_6467(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2O00F),
				.b1(W2O01F),
				.b2(W2O02F),
				.b3(W2O10F),
				.b4(W2O11F),
				.b5(W2O12F),
				.b6(W2O20F),
				.b7(W2O21F),
				.b8(W2O22F),
				.c(c2F02O)
);

assign C202O=c2002O+c2102O+c2202O+c2302O+c2402O+c2502O+c2602O+c2702O+c2802O+c2902O+c2A02O+c2B02O+c2C02O+c2D02O+c2E02O+c2F02O;
assign A202O=(C202O>=0)?1:0;

assign P302O=A202O;

ninexnine_unit ninexnine_unit_6468(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2O000),
				.b1(W2O010),
				.b2(W2O020),
				.b3(W2O100),
				.b4(W2O110),
				.b5(W2O120),
				.b6(W2O200),
				.b7(W2O210),
				.b8(W2O220),
				.c(c2010O)
);

ninexnine_unit ninexnine_unit_6469(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2O001),
				.b1(W2O011),
				.b2(W2O021),
				.b3(W2O101),
				.b4(W2O111),
				.b5(W2O121),
				.b6(W2O201),
				.b7(W2O211),
				.b8(W2O221),
				.c(c2110O)
);

ninexnine_unit ninexnine_unit_6470(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2O002),
				.b1(W2O012),
				.b2(W2O022),
				.b3(W2O102),
				.b4(W2O112),
				.b5(W2O122),
				.b6(W2O202),
				.b7(W2O212),
				.b8(W2O222),
				.c(c2210O)
);

ninexnine_unit ninexnine_unit_6471(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2O003),
				.b1(W2O013),
				.b2(W2O023),
				.b3(W2O103),
				.b4(W2O113),
				.b5(W2O123),
				.b6(W2O203),
				.b7(W2O213),
				.b8(W2O223),
				.c(c2310O)
);

ninexnine_unit ninexnine_unit_6472(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2O004),
				.b1(W2O014),
				.b2(W2O024),
				.b3(W2O104),
				.b4(W2O114),
				.b5(W2O124),
				.b6(W2O204),
				.b7(W2O214),
				.b8(W2O224),
				.c(c2410O)
);

ninexnine_unit ninexnine_unit_6473(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2O005),
				.b1(W2O015),
				.b2(W2O025),
				.b3(W2O105),
				.b4(W2O115),
				.b5(W2O125),
				.b6(W2O205),
				.b7(W2O215),
				.b8(W2O225),
				.c(c2510O)
);

ninexnine_unit ninexnine_unit_6474(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2O006),
				.b1(W2O016),
				.b2(W2O026),
				.b3(W2O106),
				.b4(W2O116),
				.b5(W2O126),
				.b6(W2O206),
				.b7(W2O216),
				.b8(W2O226),
				.c(c2610O)
);

ninexnine_unit ninexnine_unit_6475(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2O007),
				.b1(W2O017),
				.b2(W2O027),
				.b3(W2O107),
				.b4(W2O117),
				.b5(W2O127),
				.b6(W2O207),
				.b7(W2O217),
				.b8(W2O227),
				.c(c2710O)
);

ninexnine_unit ninexnine_unit_6476(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2O008),
				.b1(W2O018),
				.b2(W2O028),
				.b3(W2O108),
				.b4(W2O118),
				.b5(W2O128),
				.b6(W2O208),
				.b7(W2O218),
				.b8(W2O228),
				.c(c2810O)
);

ninexnine_unit ninexnine_unit_6477(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2O009),
				.b1(W2O019),
				.b2(W2O029),
				.b3(W2O109),
				.b4(W2O119),
				.b5(W2O129),
				.b6(W2O209),
				.b7(W2O219),
				.b8(W2O229),
				.c(c2910O)
);

ninexnine_unit ninexnine_unit_6478(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2O00A),
				.b1(W2O01A),
				.b2(W2O02A),
				.b3(W2O10A),
				.b4(W2O11A),
				.b5(W2O12A),
				.b6(W2O20A),
				.b7(W2O21A),
				.b8(W2O22A),
				.c(c2A10O)
);

ninexnine_unit ninexnine_unit_6479(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2O00B),
				.b1(W2O01B),
				.b2(W2O02B),
				.b3(W2O10B),
				.b4(W2O11B),
				.b5(W2O12B),
				.b6(W2O20B),
				.b7(W2O21B),
				.b8(W2O22B),
				.c(c2B10O)
);

ninexnine_unit ninexnine_unit_6480(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2O00C),
				.b1(W2O01C),
				.b2(W2O02C),
				.b3(W2O10C),
				.b4(W2O11C),
				.b5(W2O12C),
				.b6(W2O20C),
				.b7(W2O21C),
				.b8(W2O22C),
				.c(c2C10O)
);

ninexnine_unit ninexnine_unit_6481(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2O00D),
				.b1(W2O01D),
				.b2(W2O02D),
				.b3(W2O10D),
				.b4(W2O11D),
				.b5(W2O12D),
				.b6(W2O20D),
				.b7(W2O21D),
				.b8(W2O22D),
				.c(c2D10O)
);

ninexnine_unit ninexnine_unit_6482(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2O00E),
				.b1(W2O01E),
				.b2(W2O02E),
				.b3(W2O10E),
				.b4(W2O11E),
				.b5(W2O12E),
				.b6(W2O20E),
				.b7(W2O21E),
				.b8(W2O22E),
				.c(c2E10O)
);

ninexnine_unit ninexnine_unit_6483(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2O00F),
				.b1(W2O01F),
				.b2(W2O02F),
				.b3(W2O10F),
				.b4(W2O11F),
				.b5(W2O12F),
				.b6(W2O20F),
				.b7(W2O21F),
				.b8(W2O22F),
				.c(c2F10O)
);

assign C210O=c2010O+c2110O+c2210O+c2310O+c2410O+c2510O+c2610O+c2710O+c2810O+c2910O+c2A10O+c2B10O+c2C10O+c2D10O+c2E10O+c2F10O;
assign A210O=(C210O>=0)?1:0;

assign P310O=A210O;

ninexnine_unit ninexnine_unit_6484(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2O000),
				.b1(W2O010),
				.b2(W2O020),
				.b3(W2O100),
				.b4(W2O110),
				.b5(W2O120),
				.b6(W2O200),
				.b7(W2O210),
				.b8(W2O220),
				.c(c2011O)
);

ninexnine_unit ninexnine_unit_6485(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2O001),
				.b1(W2O011),
				.b2(W2O021),
				.b3(W2O101),
				.b4(W2O111),
				.b5(W2O121),
				.b6(W2O201),
				.b7(W2O211),
				.b8(W2O221),
				.c(c2111O)
);

ninexnine_unit ninexnine_unit_6486(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2O002),
				.b1(W2O012),
				.b2(W2O022),
				.b3(W2O102),
				.b4(W2O112),
				.b5(W2O122),
				.b6(W2O202),
				.b7(W2O212),
				.b8(W2O222),
				.c(c2211O)
);

ninexnine_unit ninexnine_unit_6487(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2O003),
				.b1(W2O013),
				.b2(W2O023),
				.b3(W2O103),
				.b4(W2O113),
				.b5(W2O123),
				.b6(W2O203),
				.b7(W2O213),
				.b8(W2O223),
				.c(c2311O)
);

ninexnine_unit ninexnine_unit_6488(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2O004),
				.b1(W2O014),
				.b2(W2O024),
				.b3(W2O104),
				.b4(W2O114),
				.b5(W2O124),
				.b6(W2O204),
				.b7(W2O214),
				.b8(W2O224),
				.c(c2411O)
);

ninexnine_unit ninexnine_unit_6489(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2O005),
				.b1(W2O015),
				.b2(W2O025),
				.b3(W2O105),
				.b4(W2O115),
				.b5(W2O125),
				.b6(W2O205),
				.b7(W2O215),
				.b8(W2O225),
				.c(c2511O)
);

ninexnine_unit ninexnine_unit_6490(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2O006),
				.b1(W2O016),
				.b2(W2O026),
				.b3(W2O106),
				.b4(W2O116),
				.b5(W2O126),
				.b6(W2O206),
				.b7(W2O216),
				.b8(W2O226),
				.c(c2611O)
);

ninexnine_unit ninexnine_unit_6491(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2O007),
				.b1(W2O017),
				.b2(W2O027),
				.b3(W2O107),
				.b4(W2O117),
				.b5(W2O127),
				.b6(W2O207),
				.b7(W2O217),
				.b8(W2O227),
				.c(c2711O)
);

ninexnine_unit ninexnine_unit_6492(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2O008),
				.b1(W2O018),
				.b2(W2O028),
				.b3(W2O108),
				.b4(W2O118),
				.b5(W2O128),
				.b6(W2O208),
				.b7(W2O218),
				.b8(W2O228),
				.c(c2811O)
);

ninexnine_unit ninexnine_unit_6493(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2O009),
				.b1(W2O019),
				.b2(W2O029),
				.b3(W2O109),
				.b4(W2O119),
				.b5(W2O129),
				.b6(W2O209),
				.b7(W2O219),
				.b8(W2O229),
				.c(c2911O)
);

ninexnine_unit ninexnine_unit_6494(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2O00A),
				.b1(W2O01A),
				.b2(W2O02A),
				.b3(W2O10A),
				.b4(W2O11A),
				.b5(W2O12A),
				.b6(W2O20A),
				.b7(W2O21A),
				.b8(W2O22A),
				.c(c2A11O)
);

ninexnine_unit ninexnine_unit_6495(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2O00B),
				.b1(W2O01B),
				.b2(W2O02B),
				.b3(W2O10B),
				.b4(W2O11B),
				.b5(W2O12B),
				.b6(W2O20B),
				.b7(W2O21B),
				.b8(W2O22B),
				.c(c2B11O)
);

ninexnine_unit ninexnine_unit_6496(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2O00C),
				.b1(W2O01C),
				.b2(W2O02C),
				.b3(W2O10C),
				.b4(W2O11C),
				.b5(W2O12C),
				.b6(W2O20C),
				.b7(W2O21C),
				.b8(W2O22C),
				.c(c2C11O)
);

ninexnine_unit ninexnine_unit_6497(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2O00D),
				.b1(W2O01D),
				.b2(W2O02D),
				.b3(W2O10D),
				.b4(W2O11D),
				.b5(W2O12D),
				.b6(W2O20D),
				.b7(W2O21D),
				.b8(W2O22D),
				.c(c2D11O)
);

ninexnine_unit ninexnine_unit_6498(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2O00E),
				.b1(W2O01E),
				.b2(W2O02E),
				.b3(W2O10E),
				.b4(W2O11E),
				.b5(W2O12E),
				.b6(W2O20E),
				.b7(W2O21E),
				.b8(W2O22E),
				.c(c2E11O)
);

ninexnine_unit ninexnine_unit_6499(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2O00F),
				.b1(W2O01F),
				.b2(W2O02F),
				.b3(W2O10F),
				.b4(W2O11F),
				.b5(W2O12F),
				.b6(W2O20F),
				.b7(W2O21F),
				.b8(W2O22F),
				.c(c2F11O)
);

assign C211O=c2011O+c2111O+c2211O+c2311O+c2411O+c2511O+c2611O+c2711O+c2811O+c2911O+c2A11O+c2B11O+c2C11O+c2D11O+c2E11O+c2F11O;
assign A211O=(C211O>=0)?1:0;

assign P311O=A211O;

ninexnine_unit ninexnine_unit_6500(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2O000),
				.b1(W2O010),
				.b2(W2O020),
				.b3(W2O100),
				.b4(W2O110),
				.b5(W2O120),
				.b6(W2O200),
				.b7(W2O210),
				.b8(W2O220),
				.c(c2012O)
);

ninexnine_unit ninexnine_unit_6501(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2O001),
				.b1(W2O011),
				.b2(W2O021),
				.b3(W2O101),
				.b4(W2O111),
				.b5(W2O121),
				.b6(W2O201),
				.b7(W2O211),
				.b8(W2O221),
				.c(c2112O)
);

ninexnine_unit ninexnine_unit_6502(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2O002),
				.b1(W2O012),
				.b2(W2O022),
				.b3(W2O102),
				.b4(W2O112),
				.b5(W2O122),
				.b6(W2O202),
				.b7(W2O212),
				.b8(W2O222),
				.c(c2212O)
);

ninexnine_unit ninexnine_unit_6503(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2O003),
				.b1(W2O013),
				.b2(W2O023),
				.b3(W2O103),
				.b4(W2O113),
				.b5(W2O123),
				.b6(W2O203),
				.b7(W2O213),
				.b8(W2O223),
				.c(c2312O)
);

ninexnine_unit ninexnine_unit_6504(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2O004),
				.b1(W2O014),
				.b2(W2O024),
				.b3(W2O104),
				.b4(W2O114),
				.b5(W2O124),
				.b6(W2O204),
				.b7(W2O214),
				.b8(W2O224),
				.c(c2412O)
);

ninexnine_unit ninexnine_unit_6505(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2O005),
				.b1(W2O015),
				.b2(W2O025),
				.b3(W2O105),
				.b4(W2O115),
				.b5(W2O125),
				.b6(W2O205),
				.b7(W2O215),
				.b8(W2O225),
				.c(c2512O)
);

ninexnine_unit ninexnine_unit_6506(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2O006),
				.b1(W2O016),
				.b2(W2O026),
				.b3(W2O106),
				.b4(W2O116),
				.b5(W2O126),
				.b6(W2O206),
				.b7(W2O216),
				.b8(W2O226),
				.c(c2612O)
);

ninexnine_unit ninexnine_unit_6507(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2O007),
				.b1(W2O017),
				.b2(W2O027),
				.b3(W2O107),
				.b4(W2O117),
				.b5(W2O127),
				.b6(W2O207),
				.b7(W2O217),
				.b8(W2O227),
				.c(c2712O)
);

ninexnine_unit ninexnine_unit_6508(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2O008),
				.b1(W2O018),
				.b2(W2O028),
				.b3(W2O108),
				.b4(W2O118),
				.b5(W2O128),
				.b6(W2O208),
				.b7(W2O218),
				.b8(W2O228),
				.c(c2812O)
);

ninexnine_unit ninexnine_unit_6509(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2O009),
				.b1(W2O019),
				.b2(W2O029),
				.b3(W2O109),
				.b4(W2O119),
				.b5(W2O129),
				.b6(W2O209),
				.b7(W2O219),
				.b8(W2O229),
				.c(c2912O)
);

ninexnine_unit ninexnine_unit_6510(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2O00A),
				.b1(W2O01A),
				.b2(W2O02A),
				.b3(W2O10A),
				.b4(W2O11A),
				.b5(W2O12A),
				.b6(W2O20A),
				.b7(W2O21A),
				.b8(W2O22A),
				.c(c2A12O)
);

ninexnine_unit ninexnine_unit_6511(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2O00B),
				.b1(W2O01B),
				.b2(W2O02B),
				.b3(W2O10B),
				.b4(W2O11B),
				.b5(W2O12B),
				.b6(W2O20B),
				.b7(W2O21B),
				.b8(W2O22B),
				.c(c2B12O)
);

ninexnine_unit ninexnine_unit_6512(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2O00C),
				.b1(W2O01C),
				.b2(W2O02C),
				.b3(W2O10C),
				.b4(W2O11C),
				.b5(W2O12C),
				.b6(W2O20C),
				.b7(W2O21C),
				.b8(W2O22C),
				.c(c2C12O)
);

ninexnine_unit ninexnine_unit_6513(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2O00D),
				.b1(W2O01D),
				.b2(W2O02D),
				.b3(W2O10D),
				.b4(W2O11D),
				.b5(W2O12D),
				.b6(W2O20D),
				.b7(W2O21D),
				.b8(W2O22D),
				.c(c2D12O)
);

ninexnine_unit ninexnine_unit_6514(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2O00E),
				.b1(W2O01E),
				.b2(W2O02E),
				.b3(W2O10E),
				.b4(W2O11E),
				.b5(W2O12E),
				.b6(W2O20E),
				.b7(W2O21E),
				.b8(W2O22E),
				.c(c2E12O)
);

ninexnine_unit ninexnine_unit_6515(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2O00F),
				.b1(W2O01F),
				.b2(W2O02F),
				.b3(W2O10F),
				.b4(W2O11F),
				.b5(W2O12F),
				.b6(W2O20F),
				.b7(W2O21F),
				.b8(W2O22F),
				.c(c2F12O)
);

assign C212O=c2012O+c2112O+c2212O+c2312O+c2412O+c2512O+c2612O+c2712O+c2812O+c2912O+c2A12O+c2B12O+c2C12O+c2D12O+c2E12O+c2F12O;
assign A212O=(C212O>=0)?1:0;

assign P312O=A212O;

ninexnine_unit ninexnine_unit_6516(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2O000),
				.b1(W2O010),
				.b2(W2O020),
				.b3(W2O100),
				.b4(W2O110),
				.b5(W2O120),
				.b6(W2O200),
				.b7(W2O210),
				.b8(W2O220),
				.c(c2020O)
);

ninexnine_unit ninexnine_unit_6517(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2O001),
				.b1(W2O011),
				.b2(W2O021),
				.b3(W2O101),
				.b4(W2O111),
				.b5(W2O121),
				.b6(W2O201),
				.b7(W2O211),
				.b8(W2O221),
				.c(c2120O)
);

ninexnine_unit ninexnine_unit_6518(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2O002),
				.b1(W2O012),
				.b2(W2O022),
				.b3(W2O102),
				.b4(W2O112),
				.b5(W2O122),
				.b6(W2O202),
				.b7(W2O212),
				.b8(W2O222),
				.c(c2220O)
);

ninexnine_unit ninexnine_unit_6519(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2O003),
				.b1(W2O013),
				.b2(W2O023),
				.b3(W2O103),
				.b4(W2O113),
				.b5(W2O123),
				.b6(W2O203),
				.b7(W2O213),
				.b8(W2O223),
				.c(c2320O)
);

ninexnine_unit ninexnine_unit_6520(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2O004),
				.b1(W2O014),
				.b2(W2O024),
				.b3(W2O104),
				.b4(W2O114),
				.b5(W2O124),
				.b6(W2O204),
				.b7(W2O214),
				.b8(W2O224),
				.c(c2420O)
);

ninexnine_unit ninexnine_unit_6521(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2O005),
				.b1(W2O015),
				.b2(W2O025),
				.b3(W2O105),
				.b4(W2O115),
				.b5(W2O125),
				.b6(W2O205),
				.b7(W2O215),
				.b8(W2O225),
				.c(c2520O)
);

ninexnine_unit ninexnine_unit_6522(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2O006),
				.b1(W2O016),
				.b2(W2O026),
				.b3(W2O106),
				.b4(W2O116),
				.b5(W2O126),
				.b6(W2O206),
				.b7(W2O216),
				.b8(W2O226),
				.c(c2620O)
);

ninexnine_unit ninexnine_unit_6523(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2O007),
				.b1(W2O017),
				.b2(W2O027),
				.b3(W2O107),
				.b4(W2O117),
				.b5(W2O127),
				.b6(W2O207),
				.b7(W2O217),
				.b8(W2O227),
				.c(c2720O)
);

ninexnine_unit ninexnine_unit_6524(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2O008),
				.b1(W2O018),
				.b2(W2O028),
				.b3(W2O108),
				.b4(W2O118),
				.b5(W2O128),
				.b6(W2O208),
				.b7(W2O218),
				.b8(W2O228),
				.c(c2820O)
);

ninexnine_unit ninexnine_unit_6525(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2O009),
				.b1(W2O019),
				.b2(W2O029),
				.b3(W2O109),
				.b4(W2O119),
				.b5(W2O129),
				.b6(W2O209),
				.b7(W2O219),
				.b8(W2O229),
				.c(c2920O)
);

ninexnine_unit ninexnine_unit_6526(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2O00A),
				.b1(W2O01A),
				.b2(W2O02A),
				.b3(W2O10A),
				.b4(W2O11A),
				.b5(W2O12A),
				.b6(W2O20A),
				.b7(W2O21A),
				.b8(W2O22A),
				.c(c2A20O)
);

ninexnine_unit ninexnine_unit_6527(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2O00B),
				.b1(W2O01B),
				.b2(W2O02B),
				.b3(W2O10B),
				.b4(W2O11B),
				.b5(W2O12B),
				.b6(W2O20B),
				.b7(W2O21B),
				.b8(W2O22B),
				.c(c2B20O)
);

ninexnine_unit ninexnine_unit_6528(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2O00C),
				.b1(W2O01C),
				.b2(W2O02C),
				.b3(W2O10C),
				.b4(W2O11C),
				.b5(W2O12C),
				.b6(W2O20C),
				.b7(W2O21C),
				.b8(W2O22C),
				.c(c2C20O)
);

ninexnine_unit ninexnine_unit_6529(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2O00D),
				.b1(W2O01D),
				.b2(W2O02D),
				.b3(W2O10D),
				.b4(W2O11D),
				.b5(W2O12D),
				.b6(W2O20D),
				.b7(W2O21D),
				.b8(W2O22D),
				.c(c2D20O)
);

ninexnine_unit ninexnine_unit_6530(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2O00E),
				.b1(W2O01E),
				.b2(W2O02E),
				.b3(W2O10E),
				.b4(W2O11E),
				.b5(W2O12E),
				.b6(W2O20E),
				.b7(W2O21E),
				.b8(W2O22E),
				.c(c2E20O)
);

ninexnine_unit ninexnine_unit_6531(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2O00F),
				.b1(W2O01F),
				.b2(W2O02F),
				.b3(W2O10F),
				.b4(W2O11F),
				.b5(W2O12F),
				.b6(W2O20F),
				.b7(W2O21F),
				.b8(W2O22F),
				.c(c2F20O)
);

assign C220O=c2020O+c2120O+c2220O+c2320O+c2420O+c2520O+c2620O+c2720O+c2820O+c2920O+c2A20O+c2B20O+c2C20O+c2D20O+c2E20O+c2F20O;
assign A220O=(C220O>=0)?1:0;

assign P320O=A220O;

ninexnine_unit ninexnine_unit_6532(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2O000),
				.b1(W2O010),
				.b2(W2O020),
				.b3(W2O100),
				.b4(W2O110),
				.b5(W2O120),
				.b6(W2O200),
				.b7(W2O210),
				.b8(W2O220),
				.c(c2021O)
);

ninexnine_unit ninexnine_unit_6533(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2O001),
				.b1(W2O011),
				.b2(W2O021),
				.b3(W2O101),
				.b4(W2O111),
				.b5(W2O121),
				.b6(W2O201),
				.b7(W2O211),
				.b8(W2O221),
				.c(c2121O)
);

ninexnine_unit ninexnine_unit_6534(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2O002),
				.b1(W2O012),
				.b2(W2O022),
				.b3(W2O102),
				.b4(W2O112),
				.b5(W2O122),
				.b6(W2O202),
				.b7(W2O212),
				.b8(W2O222),
				.c(c2221O)
);

ninexnine_unit ninexnine_unit_6535(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2O003),
				.b1(W2O013),
				.b2(W2O023),
				.b3(W2O103),
				.b4(W2O113),
				.b5(W2O123),
				.b6(W2O203),
				.b7(W2O213),
				.b8(W2O223),
				.c(c2321O)
);

ninexnine_unit ninexnine_unit_6536(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2O004),
				.b1(W2O014),
				.b2(W2O024),
				.b3(W2O104),
				.b4(W2O114),
				.b5(W2O124),
				.b6(W2O204),
				.b7(W2O214),
				.b8(W2O224),
				.c(c2421O)
);

ninexnine_unit ninexnine_unit_6537(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2O005),
				.b1(W2O015),
				.b2(W2O025),
				.b3(W2O105),
				.b4(W2O115),
				.b5(W2O125),
				.b6(W2O205),
				.b7(W2O215),
				.b8(W2O225),
				.c(c2521O)
);

ninexnine_unit ninexnine_unit_6538(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2O006),
				.b1(W2O016),
				.b2(W2O026),
				.b3(W2O106),
				.b4(W2O116),
				.b5(W2O126),
				.b6(W2O206),
				.b7(W2O216),
				.b8(W2O226),
				.c(c2621O)
);

ninexnine_unit ninexnine_unit_6539(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2O007),
				.b1(W2O017),
				.b2(W2O027),
				.b3(W2O107),
				.b4(W2O117),
				.b5(W2O127),
				.b6(W2O207),
				.b7(W2O217),
				.b8(W2O227),
				.c(c2721O)
);

ninexnine_unit ninexnine_unit_6540(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2O008),
				.b1(W2O018),
				.b2(W2O028),
				.b3(W2O108),
				.b4(W2O118),
				.b5(W2O128),
				.b6(W2O208),
				.b7(W2O218),
				.b8(W2O228),
				.c(c2821O)
);

ninexnine_unit ninexnine_unit_6541(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2O009),
				.b1(W2O019),
				.b2(W2O029),
				.b3(W2O109),
				.b4(W2O119),
				.b5(W2O129),
				.b6(W2O209),
				.b7(W2O219),
				.b8(W2O229),
				.c(c2921O)
);

ninexnine_unit ninexnine_unit_6542(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2O00A),
				.b1(W2O01A),
				.b2(W2O02A),
				.b3(W2O10A),
				.b4(W2O11A),
				.b5(W2O12A),
				.b6(W2O20A),
				.b7(W2O21A),
				.b8(W2O22A),
				.c(c2A21O)
);

ninexnine_unit ninexnine_unit_6543(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2O00B),
				.b1(W2O01B),
				.b2(W2O02B),
				.b3(W2O10B),
				.b4(W2O11B),
				.b5(W2O12B),
				.b6(W2O20B),
				.b7(W2O21B),
				.b8(W2O22B),
				.c(c2B21O)
);

ninexnine_unit ninexnine_unit_6544(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2O00C),
				.b1(W2O01C),
				.b2(W2O02C),
				.b3(W2O10C),
				.b4(W2O11C),
				.b5(W2O12C),
				.b6(W2O20C),
				.b7(W2O21C),
				.b8(W2O22C),
				.c(c2C21O)
);

ninexnine_unit ninexnine_unit_6545(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2O00D),
				.b1(W2O01D),
				.b2(W2O02D),
				.b3(W2O10D),
				.b4(W2O11D),
				.b5(W2O12D),
				.b6(W2O20D),
				.b7(W2O21D),
				.b8(W2O22D),
				.c(c2D21O)
);

ninexnine_unit ninexnine_unit_6546(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2O00E),
				.b1(W2O01E),
				.b2(W2O02E),
				.b3(W2O10E),
				.b4(W2O11E),
				.b5(W2O12E),
				.b6(W2O20E),
				.b7(W2O21E),
				.b8(W2O22E),
				.c(c2E21O)
);

ninexnine_unit ninexnine_unit_6547(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2O00F),
				.b1(W2O01F),
				.b2(W2O02F),
				.b3(W2O10F),
				.b4(W2O11F),
				.b5(W2O12F),
				.b6(W2O20F),
				.b7(W2O21F),
				.b8(W2O22F),
				.c(c2F21O)
);

assign C221O=c2021O+c2121O+c2221O+c2321O+c2421O+c2521O+c2621O+c2721O+c2821O+c2921O+c2A21O+c2B21O+c2C21O+c2D21O+c2E21O+c2F21O;
assign A221O=(C221O>=0)?1:0;

assign P321O=A221O;

ninexnine_unit ninexnine_unit_6548(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2O000),
				.b1(W2O010),
				.b2(W2O020),
				.b3(W2O100),
				.b4(W2O110),
				.b5(W2O120),
				.b6(W2O200),
				.b7(W2O210),
				.b8(W2O220),
				.c(c2022O)
);

ninexnine_unit ninexnine_unit_6549(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2O001),
				.b1(W2O011),
				.b2(W2O021),
				.b3(W2O101),
				.b4(W2O111),
				.b5(W2O121),
				.b6(W2O201),
				.b7(W2O211),
				.b8(W2O221),
				.c(c2122O)
);

ninexnine_unit ninexnine_unit_6550(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2O002),
				.b1(W2O012),
				.b2(W2O022),
				.b3(W2O102),
				.b4(W2O112),
				.b5(W2O122),
				.b6(W2O202),
				.b7(W2O212),
				.b8(W2O222),
				.c(c2222O)
);

ninexnine_unit ninexnine_unit_6551(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2O003),
				.b1(W2O013),
				.b2(W2O023),
				.b3(W2O103),
				.b4(W2O113),
				.b5(W2O123),
				.b6(W2O203),
				.b7(W2O213),
				.b8(W2O223),
				.c(c2322O)
);

ninexnine_unit ninexnine_unit_6552(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2O004),
				.b1(W2O014),
				.b2(W2O024),
				.b3(W2O104),
				.b4(W2O114),
				.b5(W2O124),
				.b6(W2O204),
				.b7(W2O214),
				.b8(W2O224),
				.c(c2422O)
);

ninexnine_unit ninexnine_unit_6553(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2O005),
				.b1(W2O015),
				.b2(W2O025),
				.b3(W2O105),
				.b4(W2O115),
				.b5(W2O125),
				.b6(W2O205),
				.b7(W2O215),
				.b8(W2O225),
				.c(c2522O)
);

ninexnine_unit ninexnine_unit_6554(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2O006),
				.b1(W2O016),
				.b2(W2O026),
				.b3(W2O106),
				.b4(W2O116),
				.b5(W2O126),
				.b6(W2O206),
				.b7(W2O216),
				.b8(W2O226),
				.c(c2622O)
);

ninexnine_unit ninexnine_unit_6555(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2O007),
				.b1(W2O017),
				.b2(W2O027),
				.b3(W2O107),
				.b4(W2O117),
				.b5(W2O127),
				.b6(W2O207),
				.b7(W2O217),
				.b8(W2O227),
				.c(c2722O)
);

ninexnine_unit ninexnine_unit_6556(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2O008),
				.b1(W2O018),
				.b2(W2O028),
				.b3(W2O108),
				.b4(W2O118),
				.b5(W2O128),
				.b6(W2O208),
				.b7(W2O218),
				.b8(W2O228),
				.c(c2822O)
);

ninexnine_unit ninexnine_unit_6557(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2O009),
				.b1(W2O019),
				.b2(W2O029),
				.b3(W2O109),
				.b4(W2O119),
				.b5(W2O129),
				.b6(W2O209),
				.b7(W2O219),
				.b8(W2O229),
				.c(c2922O)
);

ninexnine_unit ninexnine_unit_6558(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2O00A),
				.b1(W2O01A),
				.b2(W2O02A),
				.b3(W2O10A),
				.b4(W2O11A),
				.b5(W2O12A),
				.b6(W2O20A),
				.b7(W2O21A),
				.b8(W2O22A),
				.c(c2A22O)
);

ninexnine_unit ninexnine_unit_6559(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2O00B),
				.b1(W2O01B),
				.b2(W2O02B),
				.b3(W2O10B),
				.b4(W2O11B),
				.b5(W2O12B),
				.b6(W2O20B),
				.b7(W2O21B),
				.b8(W2O22B),
				.c(c2B22O)
);

ninexnine_unit ninexnine_unit_6560(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2O00C),
				.b1(W2O01C),
				.b2(W2O02C),
				.b3(W2O10C),
				.b4(W2O11C),
				.b5(W2O12C),
				.b6(W2O20C),
				.b7(W2O21C),
				.b8(W2O22C),
				.c(c2C22O)
);

ninexnine_unit ninexnine_unit_6561(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2O00D),
				.b1(W2O01D),
				.b2(W2O02D),
				.b3(W2O10D),
				.b4(W2O11D),
				.b5(W2O12D),
				.b6(W2O20D),
				.b7(W2O21D),
				.b8(W2O22D),
				.c(c2D22O)
);

ninexnine_unit ninexnine_unit_6562(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2O00E),
				.b1(W2O01E),
				.b2(W2O02E),
				.b3(W2O10E),
				.b4(W2O11E),
				.b5(W2O12E),
				.b6(W2O20E),
				.b7(W2O21E),
				.b8(W2O22E),
				.c(c2E22O)
);

ninexnine_unit ninexnine_unit_6563(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2O00F),
				.b1(W2O01F),
				.b2(W2O02F),
				.b3(W2O10F),
				.b4(W2O11F),
				.b5(W2O12F),
				.b6(W2O20F),
				.b7(W2O21F),
				.b8(W2O22F),
				.c(c2F22O)
);

assign C222O=c2022O+c2122O+c2222O+c2322O+c2422O+c2522O+c2622O+c2722O+c2822O+c2922O+c2A22O+c2B22O+c2C22O+c2D22O+c2E22O+c2F22O;
assign A222O=(C222O>=0)?1:0;

assign P322O=A222O;

ninexnine_unit ninexnine_unit_6564(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2P000),
				.b1(W2P010),
				.b2(W2P020),
				.b3(W2P100),
				.b4(W2P110),
				.b5(W2P120),
				.b6(W2P200),
				.b7(W2P210),
				.b8(W2P220),
				.c(c2000P)
);

ninexnine_unit ninexnine_unit_6565(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2P001),
				.b1(W2P011),
				.b2(W2P021),
				.b3(W2P101),
				.b4(W2P111),
				.b5(W2P121),
				.b6(W2P201),
				.b7(W2P211),
				.b8(W2P221),
				.c(c2100P)
);

ninexnine_unit ninexnine_unit_6566(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2P002),
				.b1(W2P012),
				.b2(W2P022),
				.b3(W2P102),
				.b4(W2P112),
				.b5(W2P122),
				.b6(W2P202),
				.b7(W2P212),
				.b8(W2P222),
				.c(c2200P)
);

ninexnine_unit ninexnine_unit_6567(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2P003),
				.b1(W2P013),
				.b2(W2P023),
				.b3(W2P103),
				.b4(W2P113),
				.b5(W2P123),
				.b6(W2P203),
				.b7(W2P213),
				.b8(W2P223),
				.c(c2300P)
);

ninexnine_unit ninexnine_unit_6568(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2P004),
				.b1(W2P014),
				.b2(W2P024),
				.b3(W2P104),
				.b4(W2P114),
				.b5(W2P124),
				.b6(W2P204),
				.b7(W2P214),
				.b8(W2P224),
				.c(c2400P)
);

ninexnine_unit ninexnine_unit_6569(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2P005),
				.b1(W2P015),
				.b2(W2P025),
				.b3(W2P105),
				.b4(W2P115),
				.b5(W2P125),
				.b6(W2P205),
				.b7(W2P215),
				.b8(W2P225),
				.c(c2500P)
);

ninexnine_unit ninexnine_unit_6570(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2P006),
				.b1(W2P016),
				.b2(W2P026),
				.b3(W2P106),
				.b4(W2P116),
				.b5(W2P126),
				.b6(W2P206),
				.b7(W2P216),
				.b8(W2P226),
				.c(c2600P)
);

ninexnine_unit ninexnine_unit_6571(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2P007),
				.b1(W2P017),
				.b2(W2P027),
				.b3(W2P107),
				.b4(W2P117),
				.b5(W2P127),
				.b6(W2P207),
				.b7(W2P217),
				.b8(W2P227),
				.c(c2700P)
);

ninexnine_unit ninexnine_unit_6572(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2P008),
				.b1(W2P018),
				.b2(W2P028),
				.b3(W2P108),
				.b4(W2P118),
				.b5(W2P128),
				.b6(W2P208),
				.b7(W2P218),
				.b8(W2P228),
				.c(c2800P)
);

ninexnine_unit ninexnine_unit_6573(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2P009),
				.b1(W2P019),
				.b2(W2P029),
				.b3(W2P109),
				.b4(W2P119),
				.b5(W2P129),
				.b6(W2P209),
				.b7(W2P219),
				.b8(W2P229),
				.c(c2900P)
);

ninexnine_unit ninexnine_unit_6574(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2P00A),
				.b1(W2P01A),
				.b2(W2P02A),
				.b3(W2P10A),
				.b4(W2P11A),
				.b5(W2P12A),
				.b6(W2P20A),
				.b7(W2P21A),
				.b8(W2P22A),
				.c(c2A00P)
);

ninexnine_unit ninexnine_unit_6575(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2P00B),
				.b1(W2P01B),
				.b2(W2P02B),
				.b3(W2P10B),
				.b4(W2P11B),
				.b5(W2P12B),
				.b6(W2P20B),
				.b7(W2P21B),
				.b8(W2P22B),
				.c(c2B00P)
);

ninexnine_unit ninexnine_unit_6576(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2P00C),
				.b1(W2P01C),
				.b2(W2P02C),
				.b3(W2P10C),
				.b4(W2P11C),
				.b5(W2P12C),
				.b6(W2P20C),
				.b7(W2P21C),
				.b8(W2P22C),
				.c(c2C00P)
);

ninexnine_unit ninexnine_unit_6577(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2P00D),
				.b1(W2P01D),
				.b2(W2P02D),
				.b3(W2P10D),
				.b4(W2P11D),
				.b5(W2P12D),
				.b6(W2P20D),
				.b7(W2P21D),
				.b8(W2P22D),
				.c(c2D00P)
);

ninexnine_unit ninexnine_unit_6578(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2P00E),
				.b1(W2P01E),
				.b2(W2P02E),
				.b3(W2P10E),
				.b4(W2P11E),
				.b5(W2P12E),
				.b6(W2P20E),
				.b7(W2P21E),
				.b8(W2P22E),
				.c(c2E00P)
);

ninexnine_unit ninexnine_unit_6579(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2P00F),
				.b1(W2P01F),
				.b2(W2P02F),
				.b3(W2P10F),
				.b4(W2P11F),
				.b5(W2P12F),
				.b6(W2P20F),
				.b7(W2P21F),
				.b8(W2P22F),
				.c(c2F00P)
);

assign C200P=c2000P+c2100P+c2200P+c2300P+c2400P+c2500P+c2600P+c2700P+c2800P+c2900P+c2A00P+c2B00P+c2C00P+c2D00P+c2E00P+c2F00P;
assign A200P=(C200P>=0)?1:0;

assign P300P=A200P;

ninexnine_unit ninexnine_unit_6580(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2P000),
				.b1(W2P010),
				.b2(W2P020),
				.b3(W2P100),
				.b4(W2P110),
				.b5(W2P120),
				.b6(W2P200),
				.b7(W2P210),
				.b8(W2P220),
				.c(c2001P)
);

ninexnine_unit ninexnine_unit_6581(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2P001),
				.b1(W2P011),
				.b2(W2P021),
				.b3(W2P101),
				.b4(W2P111),
				.b5(W2P121),
				.b6(W2P201),
				.b7(W2P211),
				.b8(W2P221),
				.c(c2101P)
);

ninexnine_unit ninexnine_unit_6582(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2P002),
				.b1(W2P012),
				.b2(W2P022),
				.b3(W2P102),
				.b4(W2P112),
				.b5(W2P122),
				.b6(W2P202),
				.b7(W2P212),
				.b8(W2P222),
				.c(c2201P)
);

ninexnine_unit ninexnine_unit_6583(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2P003),
				.b1(W2P013),
				.b2(W2P023),
				.b3(W2P103),
				.b4(W2P113),
				.b5(W2P123),
				.b6(W2P203),
				.b7(W2P213),
				.b8(W2P223),
				.c(c2301P)
);

ninexnine_unit ninexnine_unit_6584(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2P004),
				.b1(W2P014),
				.b2(W2P024),
				.b3(W2P104),
				.b4(W2P114),
				.b5(W2P124),
				.b6(W2P204),
				.b7(W2P214),
				.b8(W2P224),
				.c(c2401P)
);

ninexnine_unit ninexnine_unit_6585(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2P005),
				.b1(W2P015),
				.b2(W2P025),
				.b3(W2P105),
				.b4(W2P115),
				.b5(W2P125),
				.b6(W2P205),
				.b7(W2P215),
				.b8(W2P225),
				.c(c2501P)
);

ninexnine_unit ninexnine_unit_6586(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2P006),
				.b1(W2P016),
				.b2(W2P026),
				.b3(W2P106),
				.b4(W2P116),
				.b5(W2P126),
				.b6(W2P206),
				.b7(W2P216),
				.b8(W2P226),
				.c(c2601P)
);

ninexnine_unit ninexnine_unit_6587(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2P007),
				.b1(W2P017),
				.b2(W2P027),
				.b3(W2P107),
				.b4(W2P117),
				.b5(W2P127),
				.b6(W2P207),
				.b7(W2P217),
				.b8(W2P227),
				.c(c2701P)
);

ninexnine_unit ninexnine_unit_6588(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2P008),
				.b1(W2P018),
				.b2(W2P028),
				.b3(W2P108),
				.b4(W2P118),
				.b5(W2P128),
				.b6(W2P208),
				.b7(W2P218),
				.b8(W2P228),
				.c(c2801P)
);

ninexnine_unit ninexnine_unit_6589(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2P009),
				.b1(W2P019),
				.b2(W2P029),
				.b3(W2P109),
				.b4(W2P119),
				.b5(W2P129),
				.b6(W2P209),
				.b7(W2P219),
				.b8(W2P229),
				.c(c2901P)
);

ninexnine_unit ninexnine_unit_6590(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2P00A),
				.b1(W2P01A),
				.b2(W2P02A),
				.b3(W2P10A),
				.b4(W2P11A),
				.b5(W2P12A),
				.b6(W2P20A),
				.b7(W2P21A),
				.b8(W2P22A),
				.c(c2A01P)
);

ninexnine_unit ninexnine_unit_6591(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2P00B),
				.b1(W2P01B),
				.b2(W2P02B),
				.b3(W2P10B),
				.b4(W2P11B),
				.b5(W2P12B),
				.b6(W2P20B),
				.b7(W2P21B),
				.b8(W2P22B),
				.c(c2B01P)
);

ninexnine_unit ninexnine_unit_6592(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2P00C),
				.b1(W2P01C),
				.b2(W2P02C),
				.b3(W2P10C),
				.b4(W2P11C),
				.b5(W2P12C),
				.b6(W2P20C),
				.b7(W2P21C),
				.b8(W2P22C),
				.c(c2C01P)
);

ninexnine_unit ninexnine_unit_6593(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2P00D),
				.b1(W2P01D),
				.b2(W2P02D),
				.b3(W2P10D),
				.b4(W2P11D),
				.b5(W2P12D),
				.b6(W2P20D),
				.b7(W2P21D),
				.b8(W2P22D),
				.c(c2D01P)
);

ninexnine_unit ninexnine_unit_6594(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2P00E),
				.b1(W2P01E),
				.b2(W2P02E),
				.b3(W2P10E),
				.b4(W2P11E),
				.b5(W2P12E),
				.b6(W2P20E),
				.b7(W2P21E),
				.b8(W2P22E),
				.c(c2E01P)
);

ninexnine_unit ninexnine_unit_6595(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2P00F),
				.b1(W2P01F),
				.b2(W2P02F),
				.b3(W2P10F),
				.b4(W2P11F),
				.b5(W2P12F),
				.b6(W2P20F),
				.b7(W2P21F),
				.b8(W2P22F),
				.c(c2F01P)
);

assign C201P=c2001P+c2101P+c2201P+c2301P+c2401P+c2501P+c2601P+c2701P+c2801P+c2901P+c2A01P+c2B01P+c2C01P+c2D01P+c2E01P+c2F01P;
assign A201P=(C201P>=0)?1:0;

assign P301P=A201P;

ninexnine_unit ninexnine_unit_6596(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2P000),
				.b1(W2P010),
				.b2(W2P020),
				.b3(W2P100),
				.b4(W2P110),
				.b5(W2P120),
				.b6(W2P200),
				.b7(W2P210),
				.b8(W2P220),
				.c(c2002P)
);

ninexnine_unit ninexnine_unit_6597(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2P001),
				.b1(W2P011),
				.b2(W2P021),
				.b3(W2P101),
				.b4(W2P111),
				.b5(W2P121),
				.b6(W2P201),
				.b7(W2P211),
				.b8(W2P221),
				.c(c2102P)
);

ninexnine_unit ninexnine_unit_6598(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2P002),
				.b1(W2P012),
				.b2(W2P022),
				.b3(W2P102),
				.b4(W2P112),
				.b5(W2P122),
				.b6(W2P202),
				.b7(W2P212),
				.b8(W2P222),
				.c(c2202P)
);

ninexnine_unit ninexnine_unit_6599(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2P003),
				.b1(W2P013),
				.b2(W2P023),
				.b3(W2P103),
				.b4(W2P113),
				.b5(W2P123),
				.b6(W2P203),
				.b7(W2P213),
				.b8(W2P223),
				.c(c2302P)
);

ninexnine_unit ninexnine_unit_6600(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2P004),
				.b1(W2P014),
				.b2(W2P024),
				.b3(W2P104),
				.b4(W2P114),
				.b5(W2P124),
				.b6(W2P204),
				.b7(W2P214),
				.b8(W2P224),
				.c(c2402P)
);

ninexnine_unit ninexnine_unit_6601(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2P005),
				.b1(W2P015),
				.b2(W2P025),
				.b3(W2P105),
				.b4(W2P115),
				.b5(W2P125),
				.b6(W2P205),
				.b7(W2P215),
				.b8(W2P225),
				.c(c2502P)
);

ninexnine_unit ninexnine_unit_6602(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2P006),
				.b1(W2P016),
				.b2(W2P026),
				.b3(W2P106),
				.b4(W2P116),
				.b5(W2P126),
				.b6(W2P206),
				.b7(W2P216),
				.b8(W2P226),
				.c(c2602P)
);

ninexnine_unit ninexnine_unit_6603(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2P007),
				.b1(W2P017),
				.b2(W2P027),
				.b3(W2P107),
				.b4(W2P117),
				.b5(W2P127),
				.b6(W2P207),
				.b7(W2P217),
				.b8(W2P227),
				.c(c2702P)
);

ninexnine_unit ninexnine_unit_6604(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2P008),
				.b1(W2P018),
				.b2(W2P028),
				.b3(W2P108),
				.b4(W2P118),
				.b5(W2P128),
				.b6(W2P208),
				.b7(W2P218),
				.b8(W2P228),
				.c(c2802P)
);

ninexnine_unit ninexnine_unit_6605(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2P009),
				.b1(W2P019),
				.b2(W2P029),
				.b3(W2P109),
				.b4(W2P119),
				.b5(W2P129),
				.b6(W2P209),
				.b7(W2P219),
				.b8(W2P229),
				.c(c2902P)
);

ninexnine_unit ninexnine_unit_6606(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2P00A),
				.b1(W2P01A),
				.b2(W2P02A),
				.b3(W2P10A),
				.b4(W2P11A),
				.b5(W2P12A),
				.b6(W2P20A),
				.b7(W2P21A),
				.b8(W2P22A),
				.c(c2A02P)
);

ninexnine_unit ninexnine_unit_6607(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2P00B),
				.b1(W2P01B),
				.b2(W2P02B),
				.b3(W2P10B),
				.b4(W2P11B),
				.b5(W2P12B),
				.b6(W2P20B),
				.b7(W2P21B),
				.b8(W2P22B),
				.c(c2B02P)
);

ninexnine_unit ninexnine_unit_6608(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2P00C),
				.b1(W2P01C),
				.b2(W2P02C),
				.b3(W2P10C),
				.b4(W2P11C),
				.b5(W2P12C),
				.b6(W2P20C),
				.b7(W2P21C),
				.b8(W2P22C),
				.c(c2C02P)
);

ninexnine_unit ninexnine_unit_6609(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2P00D),
				.b1(W2P01D),
				.b2(W2P02D),
				.b3(W2P10D),
				.b4(W2P11D),
				.b5(W2P12D),
				.b6(W2P20D),
				.b7(W2P21D),
				.b8(W2P22D),
				.c(c2D02P)
);

ninexnine_unit ninexnine_unit_6610(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2P00E),
				.b1(W2P01E),
				.b2(W2P02E),
				.b3(W2P10E),
				.b4(W2P11E),
				.b5(W2P12E),
				.b6(W2P20E),
				.b7(W2P21E),
				.b8(W2P22E),
				.c(c2E02P)
);

ninexnine_unit ninexnine_unit_6611(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2P00F),
				.b1(W2P01F),
				.b2(W2P02F),
				.b3(W2P10F),
				.b4(W2P11F),
				.b5(W2P12F),
				.b6(W2P20F),
				.b7(W2P21F),
				.b8(W2P22F),
				.c(c2F02P)
);

assign C202P=c2002P+c2102P+c2202P+c2302P+c2402P+c2502P+c2602P+c2702P+c2802P+c2902P+c2A02P+c2B02P+c2C02P+c2D02P+c2E02P+c2F02P;
assign A202P=(C202P>=0)?1:0;

assign P302P=A202P;

ninexnine_unit ninexnine_unit_6612(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2P000),
				.b1(W2P010),
				.b2(W2P020),
				.b3(W2P100),
				.b4(W2P110),
				.b5(W2P120),
				.b6(W2P200),
				.b7(W2P210),
				.b8(W2P220),
				.c(c2010P)
);

ninexnine_unit ninexnine_unit_6613(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2P001),
				.b1(W2P011),
				.b2(W2P021),
				.b3(W2P101),
				.b4(W2P111),
				.b5(W2P121),
				.b6(W2P201),
				.b7(W2P211),
				.b8(W2P221),
				.c(c2110P)
);

ninexnine_unit ninexnine_unit_6614(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2P002),
				.b1(W2P012),
				.b2(W2P022),
				.b3(W2P102),
				.b4(W2P112),
				.b5(W2P122),
				.b6(W2P202),
				.b7(W2P212),
				.b8(W2P222),
				.c(c2210P)
);

ninexnine_unit ninexnine_unit_6615(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2P003),
				.b1(W2P013),
				.b2(W2P023),
				.b3(W2P103),
				.b4(W2P113),
				.b5(W2P123),
				.b6(W2P203),
				.b7(W2P213),
				.b8(W2P223),
				.c(c2310P)
);

ninexnine_unit ninexnine_unit_6616(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2P004),
				.b1(W2P014),
				.b2(W2P024),
				.b3(W2P104),
				.b4(W2P114),
				.b5(W2P124),
				.b6(W2P204),
				.b7(W2P214),
				.b8(W2P224),
				.c(c2410P)
);

ninexnine_unit ninexnine_unit_6617(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2P005),
				.b1(W2P015),
				.b2(W2P025),
				.b3(W2P105),
				.b4(W2P115),
				.b5(W2P125),
				.b6(W2P205),
				.b7(W2P215),
				.b8(W2P225),
				.c(c2510P)
);

ninexnine_unit ninexnine_unit_6618(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2P006),
				.b1(W2P016),
				.b2(W2P026),
				.b3(W2P106),
				.b4(W2P116),
				.b5(W2P126),
				.b6(W2P206),
				.b7(W2P216),
				.b8(W2P226),
				.c(c2610P)
);

ninexnine_unit ninexnine_unit_6619(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2P007),
				.b1(W2P017),
				.b2(W2P027),
				.b3(W2P107),
				.b4(W2P117),
				.b5(W2P127),
				.b6(W2P207),
				.b7(W2P217),
				.b8(W2P227),
				.c(c2710P)
);

ninexnine_unit ninexnine_unit_6620(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2P008),
				.b1(W2P018),
				.b2(W2P028),
				.b3(W2P108),
				.b4(W2P118),
				.b5(W2P128),
				.b6(W2P208),
				.b7(W2P218),
				.b8(W2P228),
				.c(c2810P)
);

ninexnine_unit ninexnine_unit_6621(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2P009),
				.b1(W2P019),
				.b2(W2P029),
				.b3(W2P109),
				.b4(W2P119),
				.b5(W2P129),
				.b6(W2P209),
				.b7(W2P219),
				.b8(W2P229),
				.c(c2910P)
);

ninexnine_unit ninexnine_unit_6622(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2P00A),
				.b1(W2P01A),
				.b2(W2P02A),
				.b3(W2P10A),
				.b4(W2P11A),
				.b5(W2P12A),
				.b6(W2P20A),
				.b7(W2P21A),
				.b8(W2P22A),
				.c(c2A10P)
);

ninexnine_unit ninexnine_unit_6623(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2P00B),
				.b1(W2P01B),
				.b2(W2P02B),
				.b3(W2P10B),
				.b4(W2P11B),
				.b5(W2P12B),
				.b6(W2P20B),
				.b7(W2P21B),
				.b8(W2P22B),
				.c(c2B10P)
);

ninexnine_unit ninexnine_unit_6624(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2P00C),
				.b1(W2P01C),
				.b2(W2P02C),
				.b3(W2P10C),
				.b4(W2P11C),
				.b5(W2P12C),
				.b6(W2P20C),
				.b7(W2P21C),
				.b8(W2P22C),
				.c(c2C10P)
);

ninexnine_unit ninexnine_unit_6625(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2P00D),
				.b1(W2P01D),
				.b2(W2P02D),
				.b3(W2P10D),
				.b4(W2P11D),
				.b5(W2P12D),
				.b6(W2P20D),
				.b7(W2P21D),
				.b8(W2P22D),
				.c(c2D10P)
);

ninexnine_unit ninexnine_unit_6626(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2P00E),
				.b1(W2P01E),
				.b2(W2P02E),
				.b3(W2P10E),
				.b4(W2P11E),
				.b5(W2P12E),
				.b6(W2P20E),
				.b7(W2P21E),
				.b8(W2P22E),
				.c(c2E10P)
);

ninexnine_unit ninexnine_unit_6627(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2P00F),
				.b1(W2P01F),
				.b2(W2P02F),
				.b3(W2P10F),
				.b4(W2P11F),
				.b5(W2P12F),
				.b6(W2P20F),
				.b7(W2P21F),
				.b8(W2P22F),
				.c(c2F10P)
);

assign C210P=c2010P+c2110P+c2210P+c2310P+c2410P+c2510P+c2610P+c2710P+c2810P+c2910P+c2A10P+c2B10P+c2C10P+c2D10P+c2E10P+c2F10P;
assign A210P=(C210P>=0)?1:0;

assign P310P=A210P;

ninexnine_unit ninexnine_unit_6628(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2P000),
				.b1(W2P010),
				.b2(W2P020),
				.b3(W2P100),
				.b4(W2P110),
				.b5(W2P120),
				.b6(W2P200),
				.b7(W2P210),
				.b8(W2P220),
				.c(c2011P)
);

ninexnine_unit ninexnine_unit_6629(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2P001),
				.b1(W2P011),
				.b2(W2P021),
				.b3(W2P101),
				.b4(W2P111),
				.b5(W2P121),
				.b6(W2P201),
				.b7(W2P211),
				.b8(W2P221),
				.c(c2111P)
);

ninexnine_unit ninexnine_unit_6630(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2P002),
				.b1(W2P012),
				.b2(W2P022),
				.b3(W2P102),
				.b4(W2P112),
				.b5(W2P122),
				.b6(W2P202),
				.b7(W2P212),
				.b8(W2P222),
				.c(c2211P)
);

ninexnine_unit ninexnine_unit_6631(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2P003),
				.b1(W2P013),
				.b2(W2P023),
				.b3(W2P103),
				.b4(W2P113),
				.b5(W2P123),
				.b6(W2P203),
				.b7(W2P213),
				.b8(W2P223),
				.c(c2311P)
);

ninexnine_unit ninexnine_unit_6632(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2P004),
				.b1(W2P014),
				.b2(W2P024),
				.b3(W2P104),
				.b4(W2P114),
				.b5(W2P124),
				.b6(W2P204),
				.b7(W2P214),
				.b8(W2P224),
				.c(c2411P)
);

ninexnine_unit ninexnine_unit_6633(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2P005),
				.b1(W2P015),
				.b2(W2P025),
				.b3(W2P105),
				.b4(W2P115),
				.b5(W2P125),
				.b6(W2P205),
				.b7(W2P215),
				.b8(W2P225),
				.c(c2511P)
);

ninexnine_unit ninexnine_unit_6634(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2P006),
				.b1(W2P016),
				.b2(W2P026),
				.b3(W2P106),
				.b4(W2P116),
				.b5(W2P126),
				.b6(W2P206),
				.b7(W2P216),
				.b8(W2P226),
				.c(c2611P)
);

ninexnine_unit ninexnine_unit_6635(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2P007),
				.b1(W2P017),
				.b2(W2P027),
				.b3(W2P107),
				.b4(W2P117),
				.b5(W2P127),
				.b6(W2P207),
				.b7(W2P217),
				.b8(W2P227),
				.c(c2711P)
);

ninexnine_unit ninexnine_unit_6636(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2P008),
				.b1(W2P018),
				.b2(W2P028),
				.b3(W2P108),
				.b4(W2P118),
				.b5(W2P128),
				.b6(W2P208),
				.b7(W2P218),
				.b8(W2P228),
				.c(c2811P)
);

ninexnine_unit ninexnine_unit_6637(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2P009),
				.b1(W2P019),
				.b2(W2P029),
				.b3(W2P109),
				.b4(W2P119),
				.b5(W2P129),
				.b6(W2P209),
				.b7(W2P219),
				.b8(W2P229),
				.c(c2911P)
);

ninexnine_unit ninexnine_unit_6638(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2P00A),
				.b1(W2P01A),
				.b2(W2P02A),
				.b3(W2P10A),
				.b4(W2P11A),
				.b5(W2P12A),
				.b6(W2P20A),
				.b7(W2P21A),
				.b8(W2P22A),
				.c(c2A11P)
);

ninexnine_unit ninexnine_unit_6639(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2P00B),
				.b1(W2P01B),
				.b2(W2P02B),
				.b3(W2P10B),
				.b4(W2P11B),
				.b5(W2P12B),
				.b6(W2P20B),
				.b7(W2P21B),
				.b8(W2P22B),
				.c(c2B11P)
);

ninexnine_unit ninexnine_unit_6640(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2P00C),
				.b1(W2P01C),
				.b2(W2P02C),
				.b3(W2P10C),
				.b4(W2P11C),
				.b5(W2P12C),
				.b6(W2P20C),
				.b7(W2P21C),
				.b8(W2P22C),
				.c(c2C11P)
);

ninexnine_unit ninexnine_unit_6641(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2P00D),
				.b1(W2P01D),
				.b2(W2P02D),
				.b3(W2P10D),
				.b4(W2P11D),
				.b5(W2P12D),
				.b6(W2P20D),
				.b7(W2P21D),
				.b8(W2P22D),
				.c(c2D11P)
);

ninexnine_unit ninexnine_unit_6642(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2P00E),
				.b1(W2P01E),
				.b2(W2P02E),
				.b3(W2P10E),
				.b4(W2P11E),
				.b5(W2P12E),
				.b6(W2P20E),
				.b7(W2P21E),
				.b8(W2P22E),
				.c(c2E11P)
);

ninexnine_unit ninexnine_unit_6643(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2P00F),
				.b1(W2P01F),
				.b2(W2P02F),
				.b3(W2P10F),
				.b4(W2P11F),
				.b5(W2P12F),
				.b6(W2P20F),
				.b7(W2P21F),
				.b8(W2P22F),
				.c(c2F11P)
);

assign C211P=c2011P+c2111P+c2211P+c2311P+c2411P+c2511P+c2611P+c2711P+c2811P+c2911P+c2A11P+c2B11P+c2C11P+c2D11P+c2E11P+c2F11P;
assign A211P=(C211P>=0)?1:0;

assign P311P=A211P;

ninexnine_unit ninexnine_unit_6644(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2P000),
				.b1(W2P010),
				.b2(W2P020),
				.b3(W2P100),
				.b4(W2P110),
				.b5(W2P120),
				.b6(W2P200),
				.b7(W2P210),
				.b8(W2P220),
				.c(c2012P)
);

ninexnine_unit ninexnine_unit_6645(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2P001),
				.b1(W2P011),
				.b2(W2P021),
				.b3(W2P101),
				.b4(W2P111),
				.b5(W2P121),
				.b6(W2P201),
				.b7(W2P211),
				.b8(W2P221),
				.c(c2112P)
);

ninexnine_unit ninexnine_unit_6646(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2P002),
				.b1(W2P012),
				.b2(W2P022),
				.b3(W2P102),
				.b4(W2P112),
				.b5(W2P122),
				.b6(W2P202),
				.b7(W2P212),
				.b8(W2P222),
				.c(c2212P)
);

ninexnine_unit ninexnine_unit_6647(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2P003),
				.b1(W2P013),
				.b2(W2P023),
				.b3(W2P103),
				.b4(W2P113),
				.b5(W2P123),
				.b6(W2P203),
				.b7(W2P213),
				.b8(W2P223),
				.c(c2312P)
);

ninexnine_unit ninexnine_unit_6648(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2P004),
				.b1(W2P014),
				.b2(W2P024),
				.b3(W2P104),
				.b4(W2P114),
				.b5(W2P124),
				.b6(W2P204),
				.b7(W2P214),
				.b8(W2P224),
				.c(c2412P)
);

ninexnine_unit ninexnine_unit_6649(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2P005),
				.b1(W2P015),
				.b2(W2P025),
				.b3(W2P105),
				.b4(W2P115),
				.b5(W2P125),
				.b6(W2P205),
				.b7(W2P215),
				.b8(W2P225),
				.c(c2512P)
);

ninexnine_unit ninexnine_unit_6650(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2P006),
				.b1(W2P016),
				.b2(W2P026),
				.b3(W2P106),
				.b4(W2P116),
				.b5(W2P126),
				.b6(W2P206),
				.b7(W2P216),
				.b8(W2P226),
				.c(c2612P)
);

ninexnine_unit ninexnine_unit_6651(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2P007),
				.b1(W2P017),
				.b2(W2P027),
				.b3(W2P107),
				.b4(W2P117),
				.b5(W2P127),
				.b6(W2P207),
				.b7(W2P217),
				.b8(W2P227),
				.c(c2712P)
);

ninexnine_unit ninexnine_unit_6652(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2P008),
				.b1(W2P018),
				.b2(W2P028),
				.b3(W2P108),
				.b4(W2P118),
				.b5(W2P128),
				.b6(W2P208),
				.b7(W2P218),
				.b8(W2P228),
				.c(c2812P)
);

ninexnine_unit ninexnine_unit_6653(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2P009),
				.b1(W2P019),
				.b2(W2P029),
				.b3(W2P109),
				.b4(W2P119),
				.b5(W2P129),
				.b6(W2P209),
				.b7(W2P219),
				.b8(W2P229),
				.c(c2912P)
);

ninexnine_unit ninexnine_unit_6654(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2P00A),
				.b1(W2P01A),
				.b2(W2P02A),
				.b3(W2P10A),
				.b4(W2P11A),
				.b5(W2P12A),
				.b6(W2P20A),
				.b7(W2P21A),
				.b8(W2P22A),
				.c(c2A12P)
);

ninexnine_unit ninexnine_unit_6655(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2P00B),
				.b1(W2P01B),
				.b2(W2P02B),
				.b3(W2P10B),
				.b4(W2P11B),
				.b5(W2P12B),
				.b6(W2P20B),
				.b7(W2P21B),
				.b8(W2P22B),
				.c(c2B12P)
);

ninexnine_unit ninexnine_unit_6656(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2P00C),
				.b1(W2P01C),
				.b2(W2P02C),
				.b3(W2P10C),
				.b4(W2P11C),
				.b5(W2P12C),
				.b6(W2P20C),
				.b7(W2P21C),
				.b8(W2P22C),
				.c(c2C12P)
);

ninexnine_unit ninexnine_unit_6657(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2P00D),
				.b1(W2P01D),
				.b2(W2P02D),
				.b3(W2P10D),
				.b4(W2P11D),
				.b5(W2P12D),
				.b6(W2P20D),
				.b7(W2P21D),
				.b8(W2P22D),
				.c(c2D12P)
);

ninexnine_unit ninexnine_unit_6658(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2P00E),
				.b1(W2P01E),
				.b2(W2P02E),
				.b3(W2P10E),
				.b4(W2P11E),
				.b5(W2P12E),
				.b6(W2P20E),
				.b7(W2P21E),
				.b8(W2P22E),
				.c(c2E12P)
);

ninexnine_unit ninexnine_unit_6659(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2P00F),
				.b1(W2P01F),
				.b2(W2P02F),
				.b3(W2P10F),
				.b4(W2P11F),
				.b5(W2P12F),
				.b6(W2P20F),
				.b7(W2P21F),
				.b8(W2P22F),
				.c(c2F12P)
);

assign C212P=c2012P+c2112P+c2212P+c2312P+c2412P+c2512P+c2612P+c2712P+c2812P+c2912P+c2A12P+c2B12P+c2C12P+c2D12P+c2E12P+c2F12P;
assign A212P=(C212P>=0)?1:0;

assign P312P=A212P;

ninexnine_unit ninexnine_unit_6660(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2P000),
				.b1(W2P010),
				.b2(W2P020),
				.b3(W2P100),
				.b4(W2P110),
				.b5(W2P120),
				.b6(W2P200),
				.b7(W2P210),
				.b8(W2P220),
				.c(c2020P)
);

ninexnine_unit ninexnine_unit_6661(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2P001),
				.b1(W2P011),
				.b2(W2P021),
				.b3(W2P101),
				.b4(W2P111),
				.b5(W2P121),
				.b6(W2P201),
				.b7(W2P211),
				.b8(W2P221),
				.c(c2120P)
);

ninexnine_unit ninexnine_unit_6662(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2P002),
				.b1(W2P012),
				.b2(W2P022),
				.b3(W2P102),
				.b4(W2P112),
				.b5(W2P122),
				.b6(W2P202),
				.b7(W2P212),
				.b8(W2P222),
				.c(c2220P)
);

ninexnine_unit ninexnine_unit_6663(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2P003),
				.b1(W2P013),
				.b2(W2P023),
				.b3(W2P103),
				.b4(W2P113),
				.b5(W2P123),
				.b6(W2P203),
				.b7(W2P213),
				.b8(W2P223),
				.c(c2320P)
);

ninexnine_unit ninexnine_unit_6664(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2P004),
				.b1(W2P014),
				.b2(W2P024),
				.b3(W2P104),
				.b4(W2P114),
				.b5(W2P124),
				.b6(W2P204),
				.b7(W2P214),
				.b8(W2P224),
				.c(c2420P)
);

ninexnine_unit ninexnine_unit_6665(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2P005),
				.b1(W2P015),
				.b2(W2P025),
				.b3(W2P105),
				.b4(W2P115),
				.b5(W2P125),
				.b6(W2P205),
				.b7(W2P215),
				.b8(W2P225),
				.c(c2520P)
);

ninexnine_unit ninexnine_unit_6666(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2P006),
				.b1(W2P016),
				.b2(W2P026),
				.b3(W2P106),
				.b4(W2P116),
				.b5(W2P126),
				.b6(W2P206),
				.b7(W2P216),
				.b8(W2P226),
				.c(c2620P)
);

ninexnine_unit ninexnine_unit_6667(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2P007),
				.b1(W2P017),
				.b2(W2P027),
				.b3(W2P107),
				.b4(W2P117),
				.b5(W2P127),
				.b6(W2P207),
				.b7(W2P217),
				.b8(W2P227),
				.c(c2720P)
);

ninexnine_unit ninexnine_unit_6668(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2P008),
				.b1(W2P018),
				.b2(W2P028),
				.b3(W2P108),
				.b4(W2P118),
				.b5(W2P128),
				.b6(W2P208),
				.b7(W2P218),
				.b8(W2P228),
				.c(c2820P)
);

ninexnine_unit ninexnine_unit_6669(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2P009),
				.b1(W2P019),
				.b2(W2P029),
				.b3(W2P109),
				.b4(W2P119),
				.b5(W2P129),
				.b6(W2P209),
				.b7(W2P219),
				.b8(W2P229),
				.c(c2920P)
);

ninexnine_unit ninexnine_unit_6670(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2P00A),
				.b1(W2P01A),
				.b2(W2P02A),
				.b3(W2P10A),
				.b4(W2P11A),
				.b5(W2P12A),
				.b6(W2P20A),
				.b7(W2P21A),
				.b8(W2P22A),
				.c(c2A20P)
);

ninexnine_unit ninexnine_unit_6671(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2P00B),
				.b1(W2P01B),
				.b2(W2P02B),
				.b3(W2P10B),
				.b4(W2P11B),
				.b5(W2P12B),
				.b6(W2P20B),
				.b7(W2P21B),
				.b8(W2P22B),
				.c(c2B20P)
);

ninexnine_unit ninexnine_unit_6672(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2P00C),
				.b1(W2P01C),
				.b2(W2P02C),
				.b3(W2P10C),
				.b4(W2P11C),
				.b5(W2P12C),
				.b6(W2P20C),
				.b7(W2P21C),
				.b8(W2P22C),
				.c(c2C20P)
);

ninexnine_unit ninexnine_unit_6673(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2P00D),
				.b1(W2P01D),
				.b2(W2P02D),
				.b3(W2P10D),
				.b4(W2P11D),
				.b5(W2P12D),
				.b6(W2P20D),
				.b7(W2P21D),
				.b8(W2P22D),
				.c(c2D20P)
);

ninexnine_unit ninexnine_unit_6674(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2P00E),
				.b1(W2P01E),
				.b2(W2P02E),
				.b3(W2P10E),
				.b4(W2P11E),
				.b5(W2P12E),
				.b6(W2P20E),
				.b7(W2P21E),
				.b8(W2P22E),
				.c(c2E20P)
);

ninexnine_unit ninexnine_unit_6675(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2P00F),
				.b1(W2P01F),
				.b2(W2P02F),
				.b3(W2P10F),
				.b4(W2P11F),
				.b5(W2P12F),
				.b6(W2P20F),
				.b7(W2P21F),
				.b8(W2P22F),
				.c(c2F20P)
);

assign C220P=c2020P+c2120P+c2220P+c2320P+c2420P+c2520P+c2620P+c2720P+c2820P+c2920P+c2A20P+c2B20P+c2C20P+c2D20P+c2E20P+c2F20P;
assign A220P=(C220P>=0)?1:0;

assign P320P=A220P;

ninexnine_unit ninexnine_unit_6676(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2P000),
				.b1(W2P010),
				.b2(W2P020),
				.b3(W2P100),
				.b4(W2P110),
				.b5(W2P120),
				.b6(W2P200),
				.b7(W2P210),
				.b8(W2P220),
				.c(c2021P)
);

ninexnine_unit ninexnine_unit_6677(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2P001),
				.b1(W2P011),
				.b2(W2P021),
				.b3(W2P101),
				.b4(W2P111),
				.b5(W2P121),
				.b6(W2P201),
				.b7(W2P211),
				.b8(W2P221),
				.c(c2121P)
);

ninexnine_unit ninexnine_unit_6678(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2P002),
				.b1(W2P012),
				.b2(W2P022),
				.b3(W2P102),
				.b4(W2P112),
				.b5(W2P122),
				.b6(W2P202),
				.b7(W2P212),
				.b8(W2P222),
				.c(c2221P)
);

ninexnine_unit ninexnine_unit_6679(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2P003),
				.b1(W2P013),
				.b2(W2P023),
				.b3(W2P103),
				.b4(W2P113),
				.b5(W2P123),
				.b6(W2P203),
				.b7(W2P213),
				.b8(W2P223),
				.c(c2321P)
);

ninexnine_unit ninexnine_unit_6680(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2P004),
				.b1(W2P014),
				.b2(W2P024),
				.b3(W2P104),
				.b4(W2P114),
				.b5(W2P124),
				.b6(W2P204),
				.b7(W2P214),
				.b8(W2P224),
				.c(c2421P)
);

ninexnine_unit ninexnine_unit_6681(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2P005),
				.b1(W2P015),
				.b2(W2P025),
				.b3(W2P105),
				.b4(W2P115),
				.b5(W2P125),
				.b6(W2P205),
				.b7(W2P215),
				.b8(W2P225),
				.c(c2521P)
);

ninexnine_unit ninexnine_unit_6682(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2P006),
				.b1(W2P016),
				.b2(W2P026),
				.b3(W2P106),
				.b4(W2P116),
				.b5(W2P126),
				.b6(W2P206),
				.b7(W2P216),
				.b8(W2P226),
				.c(c2621P)
);

ninexnine_unit ninexnine_unit_6683(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2P007),
				.b1(W2P017),
				.b2(W2P027),
				.b3(W2P107),
				.b4(W2P117),
				.b5(W2P127),
				.b6(W2P207),
				.b7(W2P217),
				.b8(W2P227),
				.c(c2721P)
);

ninexnine_unit ninexnine_unit_6684(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2P008),
				.b1(W2P018),
				.b2(W2P028),
				.b3(W2P108),
				.b4(W2P118),
				.b5(W2P128),
				.b6(W2P208),
				.b7(W2P218),
				.b8(W2P228),
				.c(c2821P)
);

ninexnine_unit ninexnine_unit_6685(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2P009),
				.b1(W2P019),
				.b2(W2P029),
				.b3(W2P109),
				.b4(W2P119),
				.b5(W2P129),
				.b6(W2P209),
				.b7(W2P219),
				.b8(W2P229),
				.c(c2921P)
);

ninexnine_unit ninexnine_unit_6686(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2P00A),
				.b1(W2P01A),
				.b2(W2P02A),
				.b3(W2P10A),
				.b4(W2P11A),
				.b5(W2P12A),
				.b6(W2P20A),
				.b7(W2P21A),
				.b8(W2P22A),
				.c(c2A21P)
);

ninexnine_unit ninexnine_unit_6687(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2P00B),
				.b1(W2P01B),
				.b2(W2P02B),
				.b3(W2P10B),
				.b4(W2P11B),
				.b5(W2P12B),
				.b6(W2P20B),
				.b7(W2P21B),
				.b8(W2P22B),
				.c(c2B21P)
);

ninexnine_unit ninexnine_unit_6688(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2P00C),
				.b1(W2P01C),
				.b2(W2P02C),
				.b3(W2P10C),
				.b4(W2P11C),
				.b5(W2P12C),
				.b6(W2P20C),
				.b7(W2P21C),
				.b8(W2P22C),
				.c(c2C21P)
);

ninexnine_unit ninexnine_unit_6689(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2P00D),
				.b1(W2P01D),
				.b2(W2P02D),
				.b3(W2P10D),
				.b4(W2P11D),
				.b5(W2P12D),
				.b6(W2P20D),
				.b7(W2P21D),
				.b8(W2P22D),
				.c(c2D21P)
);

ninexnine_unit ninexnine_unit_6690(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2P00E),
				.b1(W2P01E),
				.b2(W2P02E),
				.b3(W2P10E),
				.b4(W2P11E),
				.b5(W2P12E),
				.b6(W2P20E),
				.b7(W2P21E),
				.b8(W2P22E),
				.c(c2E21P)
);

ninexnine_unit ninexnine_unit_6691(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2P00F),
				.b1(W2P01F),
				.b2(W2P02F),
				.b3(W2P10F),
				.b4(W2P11F),
				.b5(W2P12F),
				.b6(W2P20F),
				.b7(W2P21F),
				.b8(W2P22F),
				.c(c2F21P)
);

assign C221P=c2021P+c2121P+c2221P+c2321P+c2421P+c2521P+c2621P+c2721P+c2821P+c2921P+c2A21P+c2B21P+c2C21P+c2D21P+c2E21P+c2F21P;
assign A221P=(C221P>=0)?1:0;

assign P321P=A221P;

ninexnine_unit ninexnine_unit_6692(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2P000),
				.b1(W2P010),
				.b2(W2P020),
				.b3(W2P100),
				.b4(W2P110),
				.b5(W2P120),
				.b6(W2P200),
				.b7(W2P210),
				.b8(W2P220),
				.c(c2022P)
);

ninexnine_unit ninexnine_unit_6693(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2P001),
				.b1(W2P011),
				.b2(W2P021),
				.b3(W2P101),
				.b4(W2P111),
				.b5(W2P121),
				.b6(W2P201),
				.b7(W2P211),
				.b8(W2P221),
				.c(c2122P)
);

ninexnine_unit ninexnine_unit_6694(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2P002),
				.b1(W2P012),
				.b2(W2P022),
				.b3(W2P102),
				.b4(W2P112),
				.b5(W2P122),
				.b6(W2P202),
				.b7(W2P212),
				.b8(W2P222),
				.c(c2222P)
);

ninexnine_unit ninexnine_unit_6695(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2P003),
				.b1(W2P013),
				.b2(W2P023),
				.b3(W2P103),
				.b4(W2P113),
				.b5(W2P123),
				.b6(W2P203),
				.b7(W2P213),
				.b8(W2P223),
				.c(c2322P)
);

ninexnine_unit ninexnine_unit_6696(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2P004),
				.b1(W2P014),
				.b2(W2P024),
				.b3(W2P104),
				.b4(W2P114),
				.b5(W2P124),
				.b6(W2P204),
				.b7(W2P214),
				.b8(W2P224),
				.c(c2422P)
);

ninexnine_unit ninexnine_unit_6697(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2P005),
				.b1(W2P015),
				.b2(W2P025),
				.b3(W2P105),
				.b4(W2P115),
				.b5(W2P125),
				.b6(W2P205),
				.b7(W2P215),
				.b8(W2P225),
				.c(c2522P)
);

ninexnine_unit ninexnine_unit_6698(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2P006),
				.b1(W2P016),
				.b2(W2P026),
				.b3(W2P106),
				.b4(W2P116),
				.b5(W2P126),
				.b6(W2P206),
				.b7(W2P216),
				.b8(W2P226),
				.c(c2622P)
);

ninexnine_unit ninexnine_unit_6699(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2P007),
				.b1(W2P017),
				.b2(W2P027),
				.b3(W2P107),
				.b4(W2P117),
				.b5(W2P127),
				.b6(W2P207),
				.b7(W2P217),
				.b8(W2P227),
				.c(c2722P)
);

ninexnine_unit ninexnine_unit_6700(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2P008),
				.b1(W2P018),
				.b2(W2P028),
				.b3(W2P108),
				.b4(W2P118),
				.b5(W2P128),
				.b6(W2P208),
				.b7(W2P218),
				.b8(W2P228),
				.c(c2822P)
);

ninexnine_unit ninexnine_unit_6701(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2P009),
				.b1(W2P019),
				.b2(W2P029),
				.b3(W2P109),
				.b4(W2P119),
				.b5(W2P129),
				.b6(W2P209),
				.b7(W2P219),
				.b8(W2P229),
				.c(c2922P)
);

ninexnine_unit ninexnine_unit_6702(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2P00A),
				.b1(W2P01A),
				.b2(W2P02A),
				.b3(W2P10A),
				.b4(W2P11A),
				.b5(W2P12A),
				.b6(W2P20A),
				.b7(W2P21A),
				.b8(W2P22A),
				.c(c2A22P)
);

ninexnine_unit ninexnine_unit_6703(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2P00B),
				.b1(W2P01B),
				.b2(W2P02B),
				.b3(W2P10B),
				.b4(W2P11B),
				.b5(W2P12B),
				.b6(W2P20B),
				.b7(W2P21B),
				.b8(W2P22B),
				.c(c2B22P)
);

ninexnine_unit ninexnine_unit_6704(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2P00C),
				.b1(W2P01C),
				.b2(W2P02C),
				.b3(W2P10C),
				.b4(W2P11C),
				.b5(W2P12C),
				.b6(W2P20C),
				.b7(W2P21C),
				.b8(W2P22C),
				.c(c2C22P)
);

ninexnine_unit ninexnine_unit_6705(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2P00D),
				.b1(W2P01D),
				.b2(W2P02D),
				.b3(W2P10D),
				.b4(W2P11D),
				.b5(W2P12D),
				.b6(W2P20D),
				.b7(W2P21D),
				.b8(W2P22D),
				.c(c2D22P)
);

ninexnine_unit ninexnine_unit_6706(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2P00E),
				.b1(W2P01E),
				.b2(W2P02E),
				.b3(W2P10E),
				.b4(W2P11E),
				.b5(W2P12E),
				.b6(W2P20E),
				.b7(W2P21E),
				.b8(W2P22E),
				.c(c2E22P)
);

ninexnine_unit ninexnine_unit_6707(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2P00F),
				.b1(W2P01F),
				.b2(W2P02F),
				.b3(W2P10F),
				.b4(W2P11F),
				.b5(W2P12F),
				.b6(W2P20F),
				.b7(W2P21F),
				.b8(W2P22F),
				.c(c2F22P)
);

assign C222P=c2022P+c2122P+c2222P+c2322P+c2422P+c2522P+c2622P+c2722P+c2822P+c2922P+c2A22P+c2B22P+c2C22P+c2D22P+c2E22P+c2F22P;
assign A222P=(C222P>=0)?1:0;

assign P322P=A222P;

ninexnine_unit ninexnine_unit_6708(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2Q000),
				.b1(W2Q010),
				.b2(W2Q020),
				.b3(W2Q100),
				.b4(W2Q110),
				.b5(W2Q120),
				.b6(W2Q200),
				.b7(W2Q210),
				.b8(W2Q220),
				.c(c2000Q)
);

ninexnine_unit ninexnine_unit_6709(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2Q001),
				.b1(W2Q011),
				.b2(W2Q021),
				.b3(W2Q101),
				.b4(W2Q111),
				.b5(W2Q121),
				.b6(W2Q201),
				.b7(W2Q211),
				.b8(W2Q221),
				.c(c2100Q)
);

ninexnine_unit ninexnine_unit_6710(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2Q002),
				.b1(W2Q012),
				.b2(W2Q022),
				.b3(W2Q102),
				.b4(W2Q112),
				.b5(W2Q122),
				.b6(W2Q202),
				.b7(W2Q212),
				.b8(W2Q222),
				.c(c2200Q)
);

ninexnine_unit ninexnine_unit_6711(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2Q003),
				.b1(W2Q013),
				.b2(W2Q023),
				.b3(W2Q103),
				.b4(W2Q113),
				.b5(W2Q123),
				.b6(W2Q203),
				.b7(W2Q213),
				.b8(W2Q223),
				.c(c2300Q)
);

ninexnine_unit ninexnine_unit_6712(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2Q004),
				.b1(W2Q014),
				.b2(W2Q024),
				.b3(W2Q104),
				.b4(W2Q114),
				.b5(W2Q124),
				.b6(W2Q204),
				.b7(W2Q214),
				.b8(W2Q224),
				.c(c2400Q)
);

ninexnine_unit ninexnine_unit_6713(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2Q005),
				.b1(W2Q015),
				.b2(W2Q025),
				.b3(W2Q105),
				.b4(W2Q115),
				.b5(W2Q125),
				.b6(W2Q205),
				.b7(W2Q215),
				.b8(W2Q225),
				.c(c2500Q)
);

ninexnine_unit ninexnine_unit_6714(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2Q006),
				.b1(W2Q016),
				.b2(W2Q026),
				.b3(W2Q106),
				.b4(W2Q116),
				.b5(W2Q126),
				.b6(W2Q206),
				.b7(W2Q216),
				.b8(W2Q226),
				.c(c2600Q)
);

ninexnine_unit ninexnine_unit_6715(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2Q007),
				.b1(W2Q017),
				.b2(W2Q027),
				.b3(W2Q107),
				.b4(W2Q117),
				.b5(W2Q127),
				.b6(W2Q207),
				.b7(W2Q217),
				.b8(W2Q227),
				.c(c2700Q)
);

ninexnine_unit ninexnine_unit_6716(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2Q008),
				.b1(W2Q018),
				.b2(W2Q028),
				.b3(W2Q108),
				.b4(W2Q118),
				.b5(W2Q128),
				.b6(W2Q208),
				.b7(W2Q218),
				.b8(W2Q228),
				.c(c2800Q)
);

ninexnine_unit ninexnine_unit_6717(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2Q009),
				.b1(W2Q019),
				.b2(W2Q029),
				.b3(W2Q109),
				.b4(W2Q119),
				.b5(W2Q129),
				.b6(W2Q209),
				.b7(W2Q219),
				.b8(W2Q229),
				.c(c2900Q)
);

ninexnine_unit ninexnine_unit_6718(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2Q00A),
				.b1(W2Q01A),
				.b2(W2Q02A),
				.b3(W2Q10A),
				.b4(W2Q11A),
				.b5(W2Q12A),
				.b6(W2Q20A),
				.b7(W2Q21A),
				.b8(W2Q22A),
				.c(c2A00Q)
);

ninexnine_unit ninexnine_unit_6719(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2Q00B),
				.b1(W2Q01B),
				.b2(W2Q02B),
				.b3(W2Q10B),
				.b4(W2Q11B),
				.b5(W2Q12B),
				.b6(W2Q20B),
				.b7(W2Q21B),
				.b8(W2Q22B),
				.c(c2B00Q)
);

ninexnine_unit ninexnine_unit_6720(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2Q00C),
				.b1(W2Q01C),
				.b2(W2Q02C),
				.b3(W2Q10C),
				.b4(W2Q11C),
				.b5(W2Q12C),
				.b6(W2Q20C),
				.b7(W2Q21C),
				.b8(W2Q22C),
				.c(c2C00Q)
);

ninexnine_unit ninexnine_unit_6721(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2Q00D),
				.b1(W2Q01D),
				.b2(W2Q02D),
				.b3(W2Q10D),
				.b4(W2Q11D),
				.b5(W2Q12D),
				.b6(W2Q20D),
				.b7(W2Q21D),
				.b8(W2Q22D),
				.c(c2D00Q)
);

ninexnine_unit ninexnine_unit_6722(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2Q00E),
				.b1(W2Q01E),
				.b2(W2Q02E),
				.b3(W2Q10E),
				.b4(W2Q11E),
				.b5(W2Q12E),
				.b6(W2Q20E),
				.b7(W2Q21E),
				.b8(W2Q22E),
				.c(c2E00Q)
);

ninexnine_unit ninexnine_unit_6723(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2Q00F),
				.b1(W2Q01F),
				.b2(W2Q02F),
				.b3(W2Q10F),
				.b4(W2Q11F),
				.b5(W2Q12F),
				.b6(W2Q20F),
				.b7(W2Q21F),
				.b8(W2Q22F),
				.c(c2F00Q)
);

assign C200Q=c2000Q+c2100Q+c2200Q+c2300Q+c2400Q+c2500Q+c2600Q+c2700Q+c2800Q+c2900Q+c2A00Q+c2B00Q+c2C00Q+c2D00Q+c2E00Q+c2F00Q;
assign A200Q=(C200Q>=0)?1:0;

assign P300Q=A200Q;

ninexnine_unit ninexnine_unit_6724(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2Q000),
				.b1(W2Q010),
				.b2(W2Q020),
				.b3(W2Q100),
				.b4(W2Q110),
				.b5(W2Q120),
				.b6(W2Q200),
				.b7(W2Q210),
				.b8(W2Q220),
				.c(c2001Q)
);

ninexnine_unit ninexnine_unit_6725(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2Q001),
				.b1(W2Q011),
				.b2(W2Q021),
				.b3(W2Q101),
				.b4(W2Q111),
				.b5(W2Q121),
				.b6(W2Q201),
				.b7(W2Q211),
				.b8(W2Q221),
				.c(c2101Q)
);

ninexnine_unit ninexnine_unit_6726(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2Q002),
				.b1(W2Q012),
				.b2(W2Q022),
				.b3(W2Q102),
				.b4(W2Q112),
				.b5(W2Q122),
				.b6(W2Q202),
				.b7(W2Q212),
				.b8(W2Q222),
				.c(c2201Q)
);

ninexnine_unit ninexnine_unit_6727(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2Q003),
				.b1(W2Q013),
				.b2(W2Q023),
				.b3(W2Q103),
				.b4(W2Q113),
				.b5(W2Q123),
				.b6(W2Q203),
				.b7(W2Q213),
				.b8(W2Q223),
				.c(c2301Q)
);

ninexnine_unit ninexnine_unit_6728(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2Q004),
				.b1(W2Q014),
				.b2(W2Q024),
				.b3(W2Q104),
				.b4(W2Q114),
				.b5(W2Q124),
				.b6(W2Q204),
				.b7(W2Q214),
				.b8(W2Q224),
				.c(c2401Q)
);

ninexnine_unit ninexnine_unit_6729(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2Q005),
				.b1(W2Q015),
				.b2(W2Q025),
				.b3(W2Q105),
				.b4(W2Q115),
				.b5(W2Q125),
				.b6(W2Q205),
				.b7(W2Q215),
				.b8(W2Q225),
				.c(c2501Q)
);

ninexnine_unit ninexnine_unit_6730(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2Q006),
				.b1(W2Q016),
				.b2(W2Q026),
				.b3(W2Q106),
				.b4(W2Q116),
				.b5(W2Q126),
				.b6(W2Q206),
				.b7(W2Q216),
				.b8(W2Q226),
				.c(c2601Q)
);

ninexnine_unit ninexnine_unit_6731(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2Q007),
				.b1(W2Q017),
				.b2(W2Q027),
				.b3(W2Q107),
				.b4(W2Q117),
				.b5(W2Q127),
				.b6(W2Q207),
				.b7(W2Q217),
				.b8(W2Q227),
				.c(c2701Q)
);

ninexnine_unit ninexnine_unit_6732(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2Q008),
				.b1(W2Q018),
				.b2(W2Q028),
				.b3(W2Q108),
				.b4(W2Q118),
				.b5(W2Q128),
				.b6(W2Q208),
				.b7(W2Q218),
				.b8(W2Q228),
				.c(c2801Q)
);

ninexnine_unit ninexnine_unit_6733(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2Q009),
				.b1(W2Q019),
				.b2(W2Q029),
				.b3(W2Q109),
				.b4(W2Q119),
				.b5(W2Q129),
				.b6(W2Q209),
				.b7(W2Q219),
				.b8(W2Q229),
				.c(c2901Q)
);

ninexnine_unit ninexnine_unit_6734(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2Q00A),
				.b1(W2Q01A),
				.b2(W2Q02A),
				.b3(W2Q10A),
				.b4(W2Q11A),
				.b5(W2Q12A),
				.b6(W2Q20A),
				.b7(W2Q21A),
				.b8(W2Q22A),
				.c(c2A01Q)
);

ninexnine_unit ninexnine_unit_6735(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2Q00B),
				.b1(W2Q01B),
				.b2(W2Q02B),
				.b3(W2Q10B),
				.b4(W2Q11B),
				.b5(W2Q12B),
				.b6(W2Q20B),
				.b7(W2Q21B),
				.b8(W2Q22B),
				.c(c2B01Q)
);

ninexnine_unit ninexnine_unit_6736(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2Q00C),
				.b1(W2Q01C),
				.b2(W2Q02C),
				.b3(W2Q10C),
				.b4(W2Q11C),
				.b5(W2Q12C),
				.b6(W2Q20C),
				.b7(W2Q21C),
				.b8(W2Q22C),
				.c(c2C01Q)
);

ninexnine_unit ninexnine_unit_6737(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2Q00D),
				.b1(W2Q01D),
				.b2(W2Q02D),
				.b3(W2Q10D),
				.b4(W2Q11D),
				.b5(W2Q12D),
				.b6(W2Q20D),
				.b7(W2Q21D),
				.b8(W2Q22D),
				.c(c2D01Q)
);

ninexnine_unit ninexnine_unit_6738(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2Q00E),
				.b1(W2Q01E),
				.b2(W2Q02E),
				.b3(W2Q10E),
				.b4(W2Q11E),
				.b5(W2Q12E),
				.b6(W2Q20E),
				.b7(W2Q21E),
				.b8(W2Q22E),
				.c(c2E01Q)
);

ninexnine_unit ninexnine_unit_6739(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2Q00F),
				.b1(W2Q01F),
				.b2(W2Q02F),
				.b3(W2Q10F),
				.b4(W2Q11F),
				.b5(W2Q12F),
				.b6(W2Q20F),
				.b7(W2Q21F),
				.b8(W2Q22F),
				.c(c2F01Q)
);

assign C201Q=c2001Q+c2101Q+c2201Q+c2301Q+c2401Q+c2501Q+c2601Q+c2701Q+c2801Q+c2901Q+c2A01Q+c2B01Q+c2C01Q+c2D01Q+c2E01Q+c2F01Q;
assign A201Q=(C201Q>=0)?1:0;

assign P301Q=A201Q;

ninexnine_unit ninexnine_unit_6740(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2Q000),
				.b1(W2Q010),
				.b2(W2Q020),
				.b3(W2Q100),
				.b4(W2Q110),
				.b5(W2Q120),
				.b6(W2Q200),
				.b7(W2Q210),
				.b8(W2Q220),
				.c(c2002Q)
);

ninexnine_unit ninexnine_unit_6741(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2Q001),
				.b1(W2Q011),
				.b2(W2Q021),
				.b3(W2Q101),
				.b4(W2Q111),
				.b5(W2Q121),
				.b6(W2Q201),
				.b7(W2Q211),
				.b8(W2Q221),
				.c(c2102Q)
);

ninexnine_unit ninexnine_unit_6742(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2Q002),
				.b1(W2Q012),
				.b2(W2Q022),
				.b3(W2Q102),
				.b4(W2Q112),
				.b5(W2Q122),
				.b6(W2Q202),
				.b7(W2Q212),
				.b8(W2Q222),
				.c(c2202Q)
);

ninexnine_unit ninexnine_unit_6743(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2Q003),
				.b1(W2Q013),
				.b2(W2Q023),
				.b3(W2Q103),
				.b4(W2Q113),
				.b5(W2Q123),
				.b6(W2Q203),
				.b7(W2Q213),
				.b8(W2Q223),
				.c(c2302Q)
);

ninexnine_unit ninexnine_unit_6744(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2Q004),
				.b1(W2Q014),
				.b2(W2Q024),
				.b3(W2Q104),
				.b4(W2Q114),
				.b5(W2Q124),
				.b6(W2Q204),
				.b7(W2Q214),
				.b8(W2Q224),
				.c(c2402Q)
);

ninexnine_unit ninexnine_unit_6745(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2Q005),
				.b1(W2Q015),
				.b2(W2Q025),
				.b3(W2Q105),
				.b4(W2Q115),
				.b5(W2Q125),
				.b6(W2Q205),
				.b7(W2Q215),
				.b8(W2Q225),
				.c(c2502Q)
);

ninexnine_unit ninexnine_unit_6746(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2Q006),
				.b1(W2Q016),
				.b2(W2Q026),
				.b3(W2Q106),
				.b4(W2Q116),
				.b5(W2Q126),
				.b6(W2Q206),
				.b7(W2Q216),
				.b8(W2Q226),
				.c(c2602Q)
);

ninexnine_unit ninexnine_unit_6747(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2Q007),
				.b1(W2Q017),
				.b2(W2Q027),
				.b3(W2Q107),
				.b4(W2Q117),
				.b5(W2Q127),
				.b6(W2Q207),
				.b7(W2Q217),
				.b8(W2Q227),
				.c(c2702Q)
);

ninexnine_unit ninexnine_unit_6748(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2Q008),
				.b1(W2Q018),
				.b2(W2Q028),
				.b3(W2Q108),
				.b4(W2Q118),
				.b5(W2Q128),
				.b6(W2Q208),
				.b7(W2Q218),
				.b8(W2Q228),
				.c(c2802Q)
);

ninexnine_unit ninexnine_unit_6749(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2Q009),
				.b1(W2Q019),
				.b2(W2Q029),
				.b3(W2Q109),
				.b4(W2Q119),
				.b5(W2Q129),
				.b6(W2Q209),
				.b7(W2Q219),
				.b8(W2Q229),
				.c(c2902Q)
);

ninexnine_unit ninexnine_unit_6750(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2Q00A),
				.b1(W2Q01A),
				.b2(W2Q02A),
				.b3(W2Q10A),
				.b4(W2Q11A),
				.b5(W2Q12A),
				.b6(W2Q20A),
				.b7(W2Q21A),
				.b8(W2Q22A),
				.c(c2A02Q)
);

ninexnine_unit ninexnine_unit_6751(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2Q00B),
				.b1(W2Q01B),
				.b2(W2Q02B),
				.b3(W2Q10B),
				.b4(W2Q11B),
				.b5(W2Q12B),
				.b6(W2Q20B),
				.b7(W2Q21B),
				.b8(W2Q22B),
				.c(c2B02Q)
);

ninexnine_unit ninexnine_unit_6752(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2Q00C),
				.b1(W2Q01C),
				.b2(W2Q02C),
				.b3(W2Q10C),
				.b4(W2Q11C),
				.b5(W2Q12C),
				.b6(W2Q20C),
				.b7(W2Q21C),
				.b8(W2Q22C),
				.c(c2C02Q)
);

ninexnine_unit ninexnine_unit_6753(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2Q00D),
				.b1(W2Q01D),
				.b2(W2Q02D),
				.b3(W2Q10D),
				.b4(W2Q11D),
				.b5(W2Q12D),
				.b6(W2Q20D),
				.b7(W2Q21D),
				.b8(W2Q22D),
				.c(c2D02Q)
);

ninexnine_unit ninexnine_unit_6754(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2Q00E),
				.b1(W2Q01E),
				.b2(W2Q02E),
				.b3(W2Q10E),
				.b4(W2Q11E),
				.b5(W2Q12E),
				.b6(W2Q20E),
				.b7(W2Q21E),
				.b8(W2Q22E),
				.c(c2E02Q)
);

ninexnine_unit ninexnine_unit_6755(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2Q00F),
				.b1(W2Q01F),
				.b2(W2Q02F),
				.b3(W2Q10F),
				.b4(W2Q11F),
				.b5(W2Q12F),
				.b6(W2Q20F),
				.b7(W2Q21F),
				.b8(W2Q22F),
				.c(c2F02Q)
);

assign C202Q=c2002Q+c2102Q+c2202Q+c2302Q+c2402Q+c2502Q+c2602Q+c2702Q+c2802Q+c2902Q+c2A02Q+c2B02Q+c2C02Q+c2D02Q+c2E02Q+c2F02Q;
assign A202Q=(C202Q>=0)?1:0;

assign P302Q=A202Q;

ninexnine_unit ninexnine_unit_6756(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2Q000),
				.b1(W2Q010),
				.b2(W2Q020),
				.b3(W2Q100),
				.b4(W2Q110),
				.b5(W2Q120),
				.b6(W2Q200),
				.b7(W2Q210),
				.b8(W2Q220),
				.c(c2010Q)
);

ninexnine_unit ninexnine_unit_6757(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2Q001),
				.b1(W2Q011),
				.b2(W2Q021),
				.b3(W2Q101),
				.b4(W2Q111),
				.b5(W2Q121),
				.b6(W2Q201),
				.b7(W2Q211),
				.b8(W2Q221),
				.c(c2110Q)
);

ninexnine_unit ninexnine_unit_6758(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2Q002),
				.b1(W2Q012),
				.b2(W2Q022),
				.b3(W2Q102),
				.b4(W2Q112),
				.b5(W2Q122),
				.b6(W2Q202),
				.b7(W2Q212),
				.b8(W2Q222),
				.c(c2210Q)
);

ninexnine_unit ninexnine_unit_6759(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2Q003),
				.b1(W2Q013),
				.b2(W2Q023),
				.b3(W2Q103),
				.b4(W2Q113),
				.b5(W2Q123),
				.b6(W2Q203),
				.b7(W2Q213),
				.b8(W2Q223),
				.c(c2310Q)
);

ninexnine_unit ninexnine_unit_6760(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2Q004),
				.b1(W2Q014),
				.b2(W2Q024),
				.b3(W2Q104),
				.b4(W2Q114),
				.b5(W2Q124),
				.b6(W2Q204),
				.b7(W2Q214),
				.b8(W2Q224),
				.c(c2410Q)
);

ninexnine_unit ninexnine_unit_6761(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2Q005),
				.b1(W2Q015),
				.b2(W2Q025),
				.b3(W2Q105),
				.b4(W2Q115),
				.b5(W2Q125),
				.b6(W2Q205),
				.b7(W2Q215),
				.b8(W2Q225),
				.c(c2510Q)
);

ninexnine_unit ninexnine_unit_6762(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2Q006),
				.b1(W2Q016),
				.b2(W2Q026),
				.b3(W2Q106),
				.b4(W2Q116),
				.b5(W2Q126),
				.b6(W2Q206),
				.b7(W2Q216),
				.b8(W2Q226),
				.c(c2610Q)
);

ninexnine_unit ninexnine_unit_6763(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2Q007),
				.b1(W2Q017),
				.b2(W2Q027),
				.b3(W2Q107),
				.b4(W2Q117),
				.b5(W2Q127),
				.b6(W2Q207),
				.b7(W2Q217),
				.b8(W2Q227),
				.c(c2710Q)
);

ninexnine_unit ninexnine_unit_6764(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2Q008),
				.b1(W2Q018),
				.b2(W2Q028),
				.b3(W2Q108),
				.b4(W2Q118),
				.b5(W2Q128),
				.b6(W2Q208),
				.b7(W2Q218),
				.b8(W2Q228),
				.c(c2810Q)
);

ninexnine_unit ninexnine_unit_6765(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2Q009),
				.b1(W2Q019),
				.b2(W2Q029),
				.b3(W2Q109),
				.b4(W2Q119),
				.b5(W2Q129),
				.b6(W2Q209),
				.b7(W2Q219),
				.b8(W2Q229),
				.c(c2910Q)
);

ninexnine_unit ninexnine_unit_6766(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2Q00A),
				.b1(W2Q01A),
				.b2(W2Q02A),
				.b3(W2Q10A),
				.b4(W2Q11A),
				.b5(W2Q12A),
				.b6(W2Q20A),
				.b7(W2Q21A),
				.b8(W2Q22A),
				.c(c2A10Q)
);

ninexnine_unit ninexnine_unit_6767(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2Q00B),
				.b1(W2Q01B),
				.b2(W2Q02B),
				.b3(W2Q10B),
				.b4(W2Q11B),
				.b5(W2Q12B),
				.b6(W2Q20B),
				.b7(W2Q21B),
				.b8(W2Q22B),
				.c(c2B10Q)
);

ninexnine_unit ninexnine_unit_6768(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2Q00C),
				.b1(W2Q01C),
				.b2(W2Q02C),
				.b3(W2Q10C),
				.b4(W2Q11C),
				.b5(W2Q12C),
				.b6(W2Q20C),
				.b7(W2Q21C),
				.b8(W2Q22C),
				.c(c2C10Q)
);

ninexnine_unit ninexnine_unit_6769(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2Q00D),
				.b1(W2Q01D),
				.b2(W2Q02D),
				.b3(W2Q10D),
				.b4(W2Q11D),
				.b5(W2Q12D),
				.b6(W2Q20D),
				.b7(W2Q21D),
				.b8(W2Q22D),
				.c(c2D10Q)
);

ninexnine_unit ninexnine_unit_6770(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2Q00E),
				.b1(W2Q01E),
				.b2(W2Q02E),
				.b3(W2Q10E),
				.b4(W2Q11E),
				.b5(W2Q12E),
				.b6(W2Q20E),
				.b7(W2Q21E),
				.b8(W2Q22E),
				.c(c2E10Q)
);

ninexnine_unit ninexnine_unit_6771(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2Q00F),
				.b1(W2Q01F),
				.b2(W2Q02F),
				.b3(W2Q10F),
				.b4(W2Q11F),
				.b5(W2Q12F),
				.b6(W2Q20F),
				.b7(W2Q21F),
				.b8(W2Q22F),
				.c(c2F10Q)
);

assign C210Q=c2010Q+c2110Q+c2210Q+c2310Q+c2410Q+c2510Q+c2610Q+c2710Q+c2810Q+c2910Q+c2A10Q+c2B10Q+c2C10Q+c2D10Q+c2E10Q+c2F10Q;
assign A210Q=(C210Q>=0)?1:0;

assign P310Q=A210Q;

ninexnine_unit ninexnine_unit_6772(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2Q000),
				.b1(W2Q010),
				.b2(W2Q020),
				.b3(W2Q100),
				.b4(W2Q110),
				.b5(W2Q120),
				.b6(W2Q200),
				.b7(W2Q210),
				.b8(W2Q220),
				.c(c2011Q)
);

ninexnine_unit ninexnine_unit_6773(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2Q001),
				.b1(W2Q011),
				.b2(W2Q021),
				.b3(W2Q101),
				.b4(W2Q111),
				.b5(W2Q121),
				.b6(W2Q201),
				.b7(W2Q211),
				.b8(W2Q221),
				.c(c2111Q)
);

ninexnine_unit ninexnine_unit_6774(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2Q002),
				.b1(W2Q012),
				.b2(W2Q022),
				.b3(W2Q102),
				.b4(W2Q112),
				.b5(W2Q122),
				.b6(W2Q202),
				.b7(W2Q212),
				.b8(W2Q222),
				.c(c2211Q)
);

ninexnine_unit ninexnine_unit_6775(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2Q003),
				.b1(W2Q013),
				.b2(W2Q023),
				.b3(W2Q103),
				.b4(W2Q113),
				.b5(W2Q123),
				.b6(W2Q203),
				.b7(W2Q213),
				.b8(W2Q223),
				.c(c2311Q)
);

ninexnine_unit ninexnine_unit_6776(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2Q004),
				.b1(W2Q014),
				.b2(W2Q024),
				.b3(W2Q104),
				.b4(W2Q114),
				.b5(W2Q124),
				.b6(W2Q204),
				.b7(W2Q214),
				.b8(W2Q224),
				.c(c2411Q)
);

ninexnine_unit ninexnine_unit_6777(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2Q005),
				.b1(W2Q015),
				.b2(W2Q025),
				.b3(W2Q105),
				.b4(W2Q115),
				.b5(W2Q125),
				.b6(W2Q205),
				.b7(W2Q215),
				.b8(W2Q225),
				.c(c2511Q)
);

ninexnine_unit ninexnine_unit_6778(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2Q006),
				.b1(W2Q016),
				.b2(W2Q026),
				.b3(W2Q106),
				.b4(W2Q116),
				.b5(W2Q126),
				.b6(W2Q206),
				.b7(W2Q216),
				.b8(W2Q226),
				.c(c2611Q)
);

ninexnine_unit ninexnine_unit_6779(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2Q007),
				.b1(W2Q017),
				.b2(W2Q027),
				.b3(W2Q107),
				.b4(W2Q117),
				.b5(W2Q127),
				.b6(W2Q207),
				.b7(W2Q217),
				.b8(W2Q227),
				.c(c2711Q)
);

ninexnine_unit ninexnine_unit_6780(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2Q008),
				.b1(W2Q018),
				.b2(W2Q028),
				.b3(W2Q108),
				.b4(W2Q118),
				.b5(W2Q128),
				.b6(W2Q208),
				.b7(W2Q218),
				.b8(W2Q228),
				.c(c2811Q)
);

ninexnine_unit ninexnine_unit_6781(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2Q009),
				.b1(W2Q019),
				.b2(W2Q029),
				.b3(W2Q109),
				.b4(W2Q119),
				.b5(W2Q129),
				.b6(W2Q209),
				.b7(W2Q219),
				.b8(W2Q229),
				.c(c2911Q)
);

ninexnine_unit ninexnine_unit_6782(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2Q00A),
				.b1(W2Q01A),
				.b2(W2Q02A),
				.b3(W2Q10A),
				.b4(W2Q11A),
				.b5(W2Q12A),
				.b6(W2Q20A),
				.b7(W2Q21A),
				.b8(W2Q22A),
				.c(c2A11Q)
);

ninexnine_unit ninexnine_unit_6783(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2Q00B),
				.b1(W2Q01B),
				.b2(W2Q02B),
				.b3(W2Q10B),
				.b4(W2Q11B),
				.b5(W2Q12B),
				.b6(W2Q20B),
				.b7(W2Q21B),
				.b8(W2Q22B),
				.c(c2B11Q)
);

ninexnine_unit ninexnine_unit_6784(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2Q00C),
				.b1(W2Q01C),
				.b2(W2Q02C),
				.b3(W2Q10C),
				.b4(W2Q11C),
				.b5(W2Q12C),
				.b6(W2Q20C),
				.b7(W2Q21C),
				.b8(W2Q22C),
				.c(c2C11Q)
);

ninexnine_unit ninexnine_unit_6785(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2Q00D),
				.b1(W2Q01D),
				.b2(W2Q02D),
				.b3(W2Q10D),
				.b4(W2Q11D),
				.b5(W2Q12D),
				.b6(W2Q20D),
				.b7(W2Q21D),
				.b8(W2Q22D),
				.c(c2D11Q)
);

ninexnine_unit ninexnine_unit_6786(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2Q00E),
				.b1(W2Q01E),
				.b2(W2Q02E),
				.b3(W2Q10E),
				.b4(W2Q11E),
				.b5(W2Q12E),
				.b6(W2Q20E),
				.b7(W2Q21E),
				.b8(W2Q22E),
				.c(c2E11Q)
);

ninexnine_unit ninexnine_unit_6787(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2Q00F),
				.b1(W2Q01F),
				.b2(W2Q02F),
				.b3(W2Q10F),
				.b4(W2Q11F),
				.b5(W2Q12F),
				.b6(W2Q20F),
				.b7(W2Q21F),
				.b8(W2Q22F),
				.c(c2F11Q)
);

assign C211Q=c2011Q+c2111Q+c2211Q+c2311Q+c2411Q+c2511Q+c2611Q+c2711Q+c2811Q+c2911Q+c2A11Q+c2B11Q+c2C11Q+c2D11Q+c2E11Q+c2F11Q;
assign A211Q=(C211Q>=0)?1:0;

assign P311Q=A211Q;

ninexnine_unit ninexnine_unit_6788(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2Q000),
				.b1(W2Q010),
				.b2(W2Q020),
				.b3(W2Q100),
				.b4(W2Q110),
				.b5(W2Q120),
				.b6(W2Q200),
				.b7(W2Q210),
				.b8(W2Q220),
				.c(c2012Q)
);

ninexnine_unit ninexnine_unit_6789(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2Q001),
				.b1(W2Q011),
				.b2(W2Q021),
				.b3(W2Q101),
				.b4(W2Q111),
				.b5(W2Q121),
				.b6(W2Q201),
				.b7(W2Q211),
				.b8(W2Q221),
				.c(c2112Q)
);

ninexnine_unit ninexnine_unit_6790(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2Q002),
				.b1(W2Q012),
				.b2(W2Q022),
				.b3(W2Q102),
				.b4(W2Q112),
				.b5(W2Q122),
				.b6(W2Q202),
				.b7(W2Q212),
				.b8(W2Q222),
				.c(c2212Q)
);

ninexnine_unit ninexnine_unit_6791(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2Q003),
				.b1(W2Q013),
				.b2(W2Q023),
				.b3(W2Q103),
				.b4(W2Q113),
				.b5(W2Q123),
				.b6(W2Q203),
				.b7(W2Q213),
				.b8(W2Q223),
				.c(c2312Q)
);

ninexnine_unit ninexnine_unit_6792(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2Q004),
				.b1(W2Q014),
				.b2(W2Q024),
				.b3(W2Q104),
				.b4(W2Q114),
				.b5(W2Q124),
				.b6(W2Q204),
				.b7(W2Q214),
				.b8(W2Q224),
				.c(c2412Q)
);

ninexnine_unit ninexnine_unit_6793(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2Q005),
				.b1(W2Q015),
				.b2(W2Q025),
				.b3(W2Q105),
				.b4(W2Q115),
				.b5(W2Q125),
				.b6(W2Q205),
				.b7(W2Q215),
				.b8(W2Q225),
				.c(c2512Q)
);

ninexnine_unit ninexnine_unit_6794(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2Q006),
				.b1(W2Q016),
				.b2(W2Q026),
				.b3(W2Q106),
				.b4(W2Q116),
				.b5(W2Q126),
				.b6(W2Q206),
				.b7(W2Q216),
				.b8(W2Q226),
				.c(c2612Q)
);

ninexnine_unit ninexnine_unit_6795(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2Q007),
				.b1(W2Q017),
				.b2(W2Q027),
				.b3(W2Q107),
				.b4(W2Q117),
				.b5(W2Q127),
				.b6(W2Q207),
				.b7(W2Q217),
				.b8(W2Q227),
				.c(c2712Q)
);

ninexnine_unit ninexnine_unit_6796(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2Q008),
				.b1(W2Q018),
				.b2(W2Q028),
				.b3(W2Q108),
				.b4(W2Q118),
				.b5(W2Q128),
				.b6(W2Q208),
				.b7(W2Q218),
				.b8(W2Q228),
				.c(c2812Q)
);

ninexnine_unit ninexnine_unit_6797(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2Q009),
				.b1(W2Q019),
				.b2(W2Q029),
				.b3(W2Q109),
				.b4(W2Q119),
				.b5(W2Q129),
				.b6(W2Q209),
				.b7(W2Q219),
				.b8(W2Q229),
				.c(c2912Q)
);

ninexnine_unit ninexnine_unit_6798(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2Q00A),
				.b1(W2Q01A),
				.b2(W2Q02A),
				.b3(W2Q10A),
				.b4(W2Q11A),
				.b5(W2Q12A),
				.b6(W2Q20A),
				.b7(W2Q21A),
				.b8(W2Q22A),
				.c(c2A12Q)
);

ninexnine_unit ninexnine_unit_6799(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2Q00B),
				.b1(W2Q01B),
				.b2(W2Q02B),
				.b3(W2Q10B),
				.b4(W2Q11B),
				.b5(W2Q12B),
				.b6(W2Q20B),
				.b7(W2Q21B),
				.b8(W2Q22B),
				.c(c2B12Q)
);

ninexnine_unit ninexnine_unit_6800(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2Q00C),
				.b1(W2Q01C),
				.b2(W2Q02C),
				.b3(W2Q10C),
				.b4(W2Q11C),
				.b5(W2Q12C),
				.b6(W2Q20C),
				.b7(W2Q21C),
				.b8(W2Q22C),
				.c(c2C12Q)
);

ninexnine_unit ninexnine_unit_6801(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2Q00D),
				.b1(W2Q01D),
				.b2(W2Q02D),
				.b3(W2Q10D),
				.b4(W2Q11D),
				.b5(W2Q12D),
				.b6(W2Q20D),
				.b7(W2Q21D),
				.b8(W2Q22D),
				.c(c2D12Q)
);

ninexnine_unit ninexnine_unit_6802(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2Q00E),
				.b1(W2Q01E),
				.b2(W2Q02E),
				.b3(W2Q10E),
				.b4(W2Q11E),
				.b5(W2Q12E),
				.b6(W2Q20E),
				.b7(W2Q21E),
				.b8(W2Q22E),
				.c(c2E12Q)
);

ninexnine_unit ninexnine_unit_6803(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2Q00F),
				.b1(W2Q01F),
				.b2(W2Q02F),
				.b3(W2Q10F),
				.b4(W2Q11F),
				.b5(W2Q12F),
				.b6(W2Q20F),
				.b7(W2Q21F),
				.b8(W2Q22F),
				.c(c2F12Q)
);

assign C212Q=c2012Q+c2112Q+c2212Q+c2312Q+c2412Q+c2512Q+c2612Q+c2712Q+c2812Q+c2912Q+c2A12Q+c2B12Q+c2C12Q+c2D12Q+c2E12Q+c2F12Q;
assign A212Q=(C212Q>=0)?1:0;

assign P312Q=A212Q;

ninexnine_unit ninexnine_unit_6804(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2Q000),
				.b1(W2Q010),
				.b2(W2Q020),
				.b3(W2Q100),
				.b4(W2Q110),
				.b5(W2Q120),
				.b6(W2Q200),
				.b7(W2Q210),
				.b8(W2Q220),
				.c(c2020Q)
);

ninexnine_unit ninexnine_unit_6805(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2Q001),
				.b1(W2Q011),
				.b2(W2Q021),
				.b3(W2Q101),
				.b4(W2Q111),
				.b5(W2Q121),
				.b6(W2Q201),
				.b7(W2Q211),
				.b8(W2Q221),
				.c(c2120Q)
);

ninexnine_unit ninexnine_unit_6806(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2Q002),
				.b1(W2Q012),
				.b2(W2Q022),
				.b3(W2Q102),
				.b4(W2Q112),
				.b5(W2Q122),
				.b6(W2Q202),
				.b7(W2Q212),
				.b8(W2Q222),
				.c(c2220Q)
);

ninexnine_unit ninexnine_unit_6807(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2Q003),
				.b1(W2Q013),
				.b2(W2Q023),
				.b3(W2Q103),
				.b4(W2Q113),
				.b5(W2Q123),
				.b6(W2Q203),
				.b7(W2Q213),
				.b8(W2Q223),
				.c(c2320Q)
);

ninexnine_unit ninexnine_unit_6808(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2Q004),
				.b1(W2Q014),
				.b2(W2Q024),
				.b3(W2Q104),
				.b4(W2Q114),
				.b5(W2Q124),
				.b6(W2Q204),
				.b7(W2Q214),
				.b8(W2Q224),
				.c(c2420Q)
);

ninexnine_unit ninexnine_unit_6809(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2Q005),
				.b1(W2Q015),
				.b2(W2Q025),
				.b3(W2Q105),
				.b4(W2Q115),
				.b5(W2Q125),
				.b6(W2Q205),
				.b7(W2Q215),
				.b8(W2Q225),
				.c(c2520Q)
);

ninexnine_unit ninexnine_unit_6810(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2Q006),
				.b1(W2Q016),
				.b2(W2Q026),
				.b3(W2Q106),
				.b4(W2Q116),
				.b5(W2Q126),
				.b6(W2Q206),
				.b7(W2Q216),
				.b8(W2Q226),
				.c(c2620Q)
);

ninexnine_unit ninexnine_unit_6811(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2Q007),
				.b1(W2Q017),
				.b2(W2Q027),
				.b3(W2Q107),
				.b4(W2Q117),
				.b5(W2Q127),
				.b6(W2Q207),
				.b7(W2Q217),
				.b8(W2Q227),
				.c(c2720Q)
);

ninexnine_unit ninexnine_unit_6812(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2Q008),
				.b1(W2Q018),
				.b2(W2Q028),
				.b3(W2Q108),
				.b4(W2Q118),
				.b5(W2Q128),
				.b6(W2Q208),
				.b7(W2Q218),
				.b8(W2Q228),
				.c(c2820Q)
);

ninexnine_unit ninexnine_unit_6813(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2Q009),
				.b1(W2Q019),
				.b2(W2Q029),
				.b3(W2Q109),
				.b4(W2Q119),
				.b5(W2Q129),
				.b6(W2Q209),
				.b7(W2Q219),
				.b8(W2Q229),
				.c(c2920Q)
);

ninexnine_unit ninexnine_unit_6814(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2Q00A),
				.b1(W2Q01A),
				.b2(W2Q02A),
				.b3(W2Q10A),
				.b4(W2Q11A),
				.b5(W2Q12A),
				.b6(W2Q20A),
				.b7(W2Q21A),
				.b8(W2Q22A),
				.c(c2A20Q)
);

ninexnine_unit ninexnine_unit_6815(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2Q00B),
				.b1(W2Q01B),
				.b2(W2Q02B),
				.b3(W2Q10B),
				.b4(W2Q11B),
				.b5(W2Q12B),
				.b6(W2Q20B),
				.b7(W2Q21B),
				.b8(W2Q22B),
				.c(c2B20Q)
);

ninexnine_unit ninexnine_unit_6816(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2Q00C),
				.b1(W2Q01C),
				.b2(W2Q02C),
				.b3(W2Q10C),
				.b4(W2Q11C),
				.b5(W2Q12C),
				.b6(W2Q20C),
				.b7(W2Q21C),
				.b8(W2Q22C),
				.c(c2C20Q)
);

ninexnine_unit ninexnine_unit_6817(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2Q00D),
				.b1(W2Q01D),
				.b2(W2Q02D),
				.b3(W2Q10D),
				.b4(W2Q11D),
				.b5(W2Q12D),
				.b6(W2Q20D),
				.b7(W2Q21D),
				.b8(W2Q22D),
				.c(c2D20Q)
);

ninexnine_unit ninexnine_unit_6818(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2Q00E),
				.b1(W2Q01E),
				.b2(W2Q02E),
				.b3(W2Q10E),
				.b4(W2Q11E),
				.b5(W2Q12E),
				.b6(W2Q20E),
				.b7(W2Q21E),
				.b8(W2Q22E),
				.c(c2E20Q)
);

ninexnine_unit ninexnine_unit_6819(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2Q00F),
				.b1(W2Q01F),
				.b2(W2Q02F),
				.b3(W2Q10F),
				.b4(W2Q11F),
				.b5(W2Q12F),
				.b6(W2Q20F),
				.b7(W2Q21F),
				.b8(W2Q22F),
				.c(c2F20Q)
);

assign C220Q=c2020Q+c2120Q+c2220Q+c2320Q+c2420Q+c2520Q+c2620Q+c2720Q+c2820Q+c2920Q+c2A20Q+c2B20Q+c2C20Q+c2D20Q+c2E20Q+c2F20Q;
assign A220Q=(C220Q>=0)?1:0;

assign P320Q=A220Q;

ninexnine_unit ninexnine_unit_6820(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2Q000),
				.b1(W2Q010),
				.b2(W2Q020),
				.b3(W2Q100),
				.b4(W2Q110),
				.b5(W2Q120),
				.b6(W2Q200),
				.b7(W2Q210),
				.b8(W2Q220),
				.c(c2021Q)
);

ninexnine_unit ninexnine_unit_6821(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2Q001),
				.b1(W2Q011),
				.b2(W2Q021),
				.b3(W2Q101),
				.b4(W2Q111),
				.b5(W2Q121),
				.b6(W2Q201),
				.b7(W2Q211),
				.b8(W2Q221),
				.c(c2121Q)
);

ninexnine_unit ninexnine_unit_6822(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2Q002),
				.b1(W2Q012),
				.b2(W2Q022),
				.b3(W2Q102),
				.b4(W2Q112),
				.b5(W2Q122),
				.b6(W2Q202),
				.b7(W2Q212),
				.b8(W2Q222),
				.c(c2221Q)
);

ninexnine_unit ninexnine_unit_6823(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2Q003),
				.b1(W2Q013),
				.b2(W2Q023),
				.b3(W2Q103),
				.b4(W2Q113),
				.b5(W2Q123),
				.b6(W2Q203),
				.b7(W2Q213),
				.b8(W2Q223),
				.c(c2321Q)
);

ninexnine_unit ninexnine_unit_6824(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2Q004),
				.b1(W2Q014),
				.b2(W2Q024),
				.b3(W2Q104),
				.b4(W2Q114),
				.b5(W2Q124),
				.b6(W2Q204),
				.b7(W2Q214),
				.b8(W2Q224),
				.c(c2421Q)
);

ninexnine_unit ninexnine_unit_6825(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2Q005),
				.b1(W2Q015),
				.b2(W2Q025),
				.b3(W2Q105),
				.b4(W2Q115),
				.b5(W2Q125),
				.b6(W2Q205),
				.b7(W2Q215),
				.b8(W2Q225),
				.c(c2521Q)
);

ninexnine_unit ninexnine_unit_6826(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2Q006),
				.b1(W2Q016),
				.b2(W2Q026),
				.b3(W2Q106),
				.b4(W2Q116),
				.b5(W2Q126),
				.b6(W2Q206),
				.b7(W2Q216),
				.b8(W2Q226),
				.c(c2621Q)
);

ninexnine_unit ninexnine_unit_6827(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2Q007),
				.b1(W2Q017),
				.b2(W2Q027),
				.b3(W2Q107),
				.b4(W2Q117),
				.b5(W2Q127),
				.b6(W2Q207),
				.b7(W2Q217),
				.b8(W2Q227),
				.c(c2721Q)
);

ninexnine_unit ninexnine_unit_6828(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2Q008),
				.b1(W2Q018),
				.b2(W2Q028),
				.b3(W2Q108),
				.b4(W2Q118),
				.b5(W2Q128),
				.b6(W2Q208),
				.b7(W2Q218),
				.b8(W2Q228),
				.c(c2821Q)
);

ninexnine_unit ninexnine_unit_6829(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2Q009),
				.b1(W2Q019),
				.b2(W2Q029),
				.b3(W2Q109),
				.b4(W2Q119),
				.b5(W2Q129),
				.b6(W2Q209),
				.b7(W2Q219),
				.b8(W2Q229),
				.c(c2921Q)
);

ninexnine_unit ninexnine_unit_6830(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2Q00A),
				.b1(W2Q01A),
				.b2(W2Q02A),
				.b3(W2Q10A),
				.b4(W2Q11A),
				.b5(W2Q12A),
				.b6(W2Q20A),
				.b7(W2Q21A),
				.b8(W2Q22A),
				.c(c2A21Q)
);

ninexnine_unit ninexnine_unit_6831(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2Q00B),
				.b1(W2Q01B),
				.b2(W2Q02B),
				.b3(W2Q10B),
				.b4(W2Q11B),
				.b5(W2Q12B),
				.b6(W2Q20B),
				.b7(W2Q21B),
				.b8(W2Q22B),
				.c(c2B21Q)
);

ninexnine_unit ninexnine_unit_6832(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2Q00C),
				.b1(W2Q01C),
				.b2(W2Q02C),
				.b3(W2Q10C),
				.b4(W2Q11C),
				.b5(W2Q12C),
				.b6(W2Q20C),
				.b7(W2Q21C),
				.b8(W2Q22C),
				.c(c2C21Q)
);

ninexnine_unit ninexnine_unit_6833(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2Q00D),
				.b1(W2Q01D),
				.b2(W2Q02D),
				.b3(W2Q10D),
				.b4(W2Q11D),
				.b5(W2Q12D),
				.b6(W2Q20D),
				.b7(W2Q21D),
				.b8(W2Q22D),
				.c(c2D21Q)
);

ninexnine_unit ninexnine_unit_6834(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2Q00E),
				.b1(W2Q01E),
				.b2(W2Q02E),
				.b3(W2Q10E),
				.b4(W2Q11E),
				.b5(W2Q12E),
				.b6(W2Q20E),
				.b7(W2Q21E),
				.b8(W2Q22E),
				.c(c2E21Q)
);

ninexnine_unit ninexnine_unit_6835(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2Q00F),
				.b1(W2Q01F),
				.b2(W2Q02F),
				.b3(W2Q10F),
				.b4(W2Q11F),
				.b5(W2Q12F),
				.b6(W2Q20F),
				.b7(W2Q21F),
				.b8(W2Q22F),
				.c(c2F21Q)
);

assign C221Q=c2021Q+c2121Q+c2221Q+c2321Q+c2421Q+c2521Q+c2621Q+c2721Q+c2821Q+c2921Q+c2A21Q+c2B21Q+c2C21Q+c2D21Q+c2E21Q+c2F21Q;
assign A221Q=(C221Q>=0)?1:0;

assign P321Q=A221Q;

ninexnine_unit ninexnine_unit_6836(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2Q000),
				.b1(W2Q010),
				.b2(W2Q020),
				.b3(W2Q100),
				.b4(W2Q110),
				.b5(W2Q120),
				.b6(W2Q200),
				.b7(W2Q210),
				.b8(W2Q220),
				.c(c2022Q)
);

ninexnine_unit ninexnine_unit_6837(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2Q001),
				.b1(W2Q011),
				.b2(W2Q021),
				.b3(W2Q101),
				.b4(W2Q111),
				.b5(W2Q121),
				.b6(W2Q201),
				.b7(W2Q211),
				.b8(W2Q221),
				.c(c2122Q)
);

ninexnine_unit ninexnine_unit_6838(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2Q002),
				.b1(W2Q012),
				.b2(W2Q022),
				.b3(W2Q102),
				.b4(W2Q112),
				.b5(W2Q122),
				.b6(W2Q202),
				.b7(W2Q212),
				.b8(W2Q222),
				.c(c2222Q)
);

ninexnine_unit ninexnine_unit_6839(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2Q003),
				.b1(W2Q013),
				.b2(W2Q023),
				.b3(W2Q103),
				.b4(W2Q113),
				.b5(W2Q123),
				.b6(W2Q203),
				.b7(W2Q213),
				.b8(W2Q223),
				.c(c2322Q)
);

ninexnine_unit ninexnine_unit_6840(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2Q004),
				.b1(W2Q014),
				.b2(W2Q024),
				.b3(W2Q104),
				.b4(W2Q114),
				.b5(W2Q124),
				.b6(W2Q204),
				.b7(W2Q214),
				.b8(W2Q224),
				.c(c2422Q)
);

ninexnine_unit ninexnine_unit_6841(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2Q005),
				.b1(W2Q015),
				.b2(W2Q025),
				.b3(W2Q105),
				.b4(W2Q115),
				.b5(W2Q125),
				.b6(W2Q205),
				.b7(W2Q215),
				.b8(W2Q225),
				.c(c2522Q)
);

ninexnine_unit ninexnine_unit_6842(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2Q006),
				.b1(W2Q016),
				.b2(W2Q026),
				.b3(W2Q106),
				.b4(W2Q116),
				.b5(W2Q126),
				.b6(W2Q206),
				.b7(W2Q216),
				.b8(W2Q226),
				.c(c2622Q)
);

ninexnine_unit ninexnine_unit_6843(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2Q007),
				.b1(W2Q017),
				.b2(W2Q027),
				.b3(W2Q107),
				.b4(W2Q117),
				.b5(W2Q127),
				.b6(W2Q207),
				.b7(W2Q217),
				.b8(W2Q227),
				.c(c2722Q)
);

ninexnine_unit ninexnine_unit_6844(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2Q008),
				.b1(W2Q018),
				.b2(W2Q028),
				.b3(W2Q108),
				.b4(W2Q118),
				.b5(W2Q128),
				.b6(W2Q208),
				.b7(W2Q218),
				.b8(W2Q228),
				.c(c2822Q)
);

ninexnine_unit ninexnine_unit_6845(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2Q009),
				.b1(W2Q019),
				.b2(W2Q029),
				.b3(W2Q109),
				.b4(W2Q119),
				.b5(W2Q129),
				.b6(W2Q209),
				.b7(W2Q219),
				.b8(W2Q229),
				.c(c2922Q)
);

ninexnine_unit ninexnine_unit_6846(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2Q00A),
				.b1(W2Q01A),
				.b2(W2Q02A),
				.b3(W2Q10A),
				.b4(W2Q11A),
				.b5(W2Q12A),
				.b6(W2Q20A),
				.b7(W2Q21A),
				.b8(W2Q22A),
				.c(c2A22Q)
);

ninexnine_unit ninexnine_unit_6847(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2Q00B),
				.b1(W2Q01B),
				.b2(W2Q02B),
				.b3(W2Q10B),
				.b4(W2Q11B),
				.b5(W2Q12B),
				.b6(W2Q20B),
				.b7(W2Q21B),
				.b8(W2Q22B),
				.c(c2B22Q)
);

ninexnine_unit ninexnine_unit_6848(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2Q00C),
				.b1(W2Q01C),
				.b2(W2Q02C),
				.b3(W2Q10C),
				.b4(W2Q11C),
				.b5(W2Q12C),
				.b6(W2Q20C),
				.b7(W2Q21C),
				.b8(W2Q22C),
				.c(c2C22Q)
);

ninexnine_unit ninexnine_unit_6849(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2Q00D),
				.b1(W2Q01D),
				.b2(W2Q02D),
				.b3(W2Q10D),
				.b4(W2Q11D),
				.b5(W2Q12D),
				.b6(W2Q20D),
				.b7(W2Q21D),
				.b8(W2Q22D),
				.c(c2D22Q)
);

ninexnine_unit ninexnine_unit_6850(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2Q00E),
				.b1(W2Q01E),
				.b2(W2Q02E),
				.b3(W2Q10E),
				.b4(W2Q11E),
				.b5(W2Q12E),
				.b6(W2Q20E),
				.b7(W2Q21E),
				.b8(W2Q22E),
				.c(c2E22Q)
);

ninexnine_unit ninexnine_unit_6851(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2Q00F),
				.b1(W2Q01F),
				.b2(W2Q02F),
				.b3(W2Q10F),
				.b4(W2Q11F),
				.b5(W2Q12F),
				.b6(W2Q20F),
				.b7(W2Q21F),
				.b8(W2Q22F),
				.c(c2F22Q)
);

assign C222Q=c2022Q+c2122Q+c2222Q+c2322Q+c2422Q+c2522Q+c2622Q+c2722Q+c2822Q+c2922Q+c2A22Q+c2B22Q+c2C22Q+c2D22Q+c2E22Q+c2F22Q;
assign A222Q=(C222Q>=0)?1:0;

assign P322Q=A222Q;

ninexnine_unit ninexnine_unit_6852(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2R000),
				.b1(W2R010),
				.b2(W2R020),
				.b3(W2R100),
				.b4(W2R110),
				.b5(W2R120),
				.b6(W2R200),
				.b7(W2R210),
				.b8(W2R220),
				.c(c2000R)
);

ninexnine_unit ninexnine_unit_6853(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2R001),
				.b1(W2R011),
				.b2(W2R021),
				.b3(W2R101),
				.b4(W2R111),
				.b5(W2R121),
				.b6(W2R201),
				.b7(W2R211),
				.b8(W2R221),
				.c(c2100R)
);

ninexnine_unit ninexnine_unit_6854(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2R002),
				.b1(W2R012),
				.b2(W2R022),
				.b3(W2R102),
				.b4(W2R112),
				.b5(W2R122),
				.b6(W2R202),
				.b7(W2R212),
				.b8(W2R222),
				.c(c2200R)
);

ninexnine_unit ninexnine_unit_6855(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2R003),
				.b1(W2R013),
				.b2(W2R023),
				.b3(W2R103),
				.b4(W2R113),
				.b5(W2R123),
				.b6(W2R203),
				.b7(W2R213),
				.b8(W2R223),
				.c(c2300R)
);

ninexnine_unit ninexnine_unit_6856(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2R004),
				.b1(W2R014),
				.b2(W2R024),
				.b3(W2R104),
				.b4(W2R114),
				.b5(W2R124),
				.b6(W2R204),
				.b7(W2R214),
				.b8(W2R224),
				.c(c2400R)
);

ninexnine_unit ninexnine_unit_6857(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2R005),
				.b1(W2R015),
				.b2(W2R025),
				.b3(W2R105),
				.b4(W2R115),
				.b5(W2R125),
				.b6(W2R205),
				.b7(W2R215),
				.b8(W2R225),
				.c(c2500R)
);

ninexnine_unit ninexnine_unit_6858(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2R006),
				.b1(W2R016),
				.b2(W2R026),
				.b3(W2R106),
				.b4(W2R116),
				.b5(W2R126),
				.b6(W2R206),
				.b7(W2R216),
				.b8(W2R226),
				.c(c2600R)
);

ninexnine_unit ninexnine_unit_6859(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2R007),
				.b1(W2R017),
				.b2(W2R027),
				.b3(W2R107),
				.b4(W2R117),
				.b5(W2R127),
				.b6(W2R207),
				.b7(W2R217),
				.b8(W2R227),
				.c(c2700R)
);

ninexnine_unit ninexnine_unit_6860(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2R008),
				.b1(W2R018),
				.b2(W2R028),
				.b3(W2R108),
				.b4(W2R118),
				.b5(W2R128),
				.b6(W2R208),
				.b7(W2R218),
				.b8(W2R228),
				.c(c2800R)
);

ninexnine_unit ninexnine_unit_6861(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2R009),
				.b1(W2R019),
				.b2(W2R029),
				.b3(W2R109),
				.b4(W2R119),
				.b5(W2R129),
				.b6(W2R209),
				.b7(W2R219),
				.b8(W2R229),
				.c(c2900R)
);

ninexnine_unit ninexnine_unit_6862(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2R00A),
				.b1(W2R01A),
				.b2(W2R02A),
				.b3(W2R10A),
				.b4(W2R11A),
				.b5(W2R12A),
				.b6(W2R20A),
				.b7(W2R21A),
				.b8(W2R22A),
				.c(c2A00R)
);

ninexnine_unit ninexnine_unit_6863(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2R00B),
				.b1(W2R01B),
				.b2(W2R02B),
				.b3(W2R10B),
				.b4(W2R11B),
				.b5(W2R12B),
				.b6(W2R20B),
				.b7(W2R21B),
				.b8(W2R22B),
				.c(c2B00R)
);

ninexnine_unit ninexnine_unit_6864(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2R00C),
				.b1(W2R01C),
				.b2(W2R02C),
				.b3(W2R10C),
				.b4(W2R11C),
				.b5(W2R12C),
				.b6(W2R20C),
				.b7(W2R21C),
				.b8(W2R22C),
				.c(c2C00R)
);

ninexnine_unit ninexnine_unit_6865(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2R00D),
				.b1(W2R01D),
				.b2(W2R02D),
				.b3(W2R10D),
				.b4(W2R11D),
				.b5(W2R12D),
				.b6(W2R20D),
				.b7(W2R21D),
				.b8(W2R22D),
				.c(c2D00R)
);

ninexnine_unit ninexnine_unit_6866(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2R00E),
				.b1(W2R01E),
				.b2(W2R02E),
				.b3(W2R10E),
				.b4(W2R11E),
				.b5(W2R12E),
				.b6(W2R20E),
				.b7(W2R21E),
				.b8(W2R22E),
				.c(c2E00R)
);

ninexnine_unit ninexnine_unit_6867(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2R00F),
				.b1(W2R01F),
				.b2(W2R02F),
				.b3(W2R10F),
				.b4(W2R11F),
				.b5(W2R12F),
				.b6(W2R20F),
				.b7(W2R21F),
				.b8(W2R22F),
				.c(c2F00R)
);

assign C200R=c2000R+c2100R+c2200R+c2300R+c2400R+c2500R+c2600R+c2700R+c2800R+c2900R+c2A00R+c2B00R+c2C00R+c2D00R+c2E00R+c2F00R;
assign A200R=(C200R>=0)?1:0;

assign P300R=A200R;

ninexnine_unit ninexnine_unit_6868(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2R000),
				.b1(W2R010),
				.b2(W2R020),
				.b3(W2R100),
				.b4(W2R110),
				.b5(W2R120),
				.b6(W2R200),
				.b7(W2R210),
				.b8(W2R220),
				.c(c2001R)
);

ninexnine_unit ninexnine_unit_6869(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2R001),
				.b1(W2R011),
				.b2(W2R021),
				.b3(W2R101),
				.b4(W2R111),
				.b5(W2R121),
				.b6(W2R201),
				.b7(W2R211),
				.b8(W2R221),
				.c(c2101R)
);

ninexnine_unit ninexnine_unit_6870(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2R002),
				.b1(W2R012),
				.b2(W2R022),
				.b3(W2R102),
				.b4(W2R112),
				.b5(W2R122),
				.b6(W2R202),
				.b7(W2R212),
				.b8(W2R222),
				.c(c2201R)
);

ninexnine_unit ninexnine_unit_6871(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2R003),
				.b1(W2R013),
				.b2(W2R023),
				.b3(W2R103),
				.b4(W2R113),
				.b5(W2R123),
				.b6(W2R203),
				.b7(W2R213),
				.b8(W2R223),
				.c(c2301R)
);

ninexnine_unit ninexnine_unit_6872(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2R004),
				.b1(W2R014),
				.b2(W2R024),
				.b3(W2R104),
				.b4(W2R114),
				.b5(W2R124),
				.b6(W2R204),
				.b7(W2R214),
				.b8(W2R224),
				.c(c2401R)
);

ninexnine_unit ninexnine_unit_6873(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2R005),
				.b1(W2R015),
				.b2(W2R025),
				.b3(W2R105),
				.b4(W2R115),
				.b5(W2R125),
				.b6(W2R205),
				.b7(W2R215),
				.b8(W2R225),
				.c(c2501R)
);

ninexnine_unit ninexnine_unit_6874(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2R006),
				.b1(W2R016),
				.b2(W2R026),
				.b3(W2R106),
				.b4(W2R116),
				.b5(W2R126),
				.b6(W2R206),
				.b7(W2R216),
				.b8(W2R226),
				.c(c2601R)
);

ninexnine_unit ninexnine_unit_6875(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2R007),
				.b1(W2R017),
				.b2(W2R027),
				.b3(W2R107),
				.b4(W2R117),
				.b5(W2R127),
				.b6(W2R207),
				.b7(W2R217),
				.b8(W2R227),
				.c(c2701R)
);

ninexnine_unit ninexnine_unit_6876(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2R008),
				.b1(W2R018),
				.b2(W2R028),
				.b3(W2R108),
				.b4(W2R118),
				.b5(W2R128),
				.b6(W2R208),
				.b7(W2R218),
				.b8(W2R228),
				.c(c2801R)
);

ninexnine_unit ninexnine_unit_6877(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2R009),
				.b1(W2R019),
				.b2(W2R029),
				.b3(W2R109),
				.b4(W2R119),
				.b5(W2R129),
				.b6(W2R209),
				.b7(W2R219),
				.b8(W2R229),
				.c(c2901R)
);

ninexnine_unit ninexnine_unit_6878(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2R00A),
				.b1(W2R01A),
				.b2(W2R02A),
				.b3(W2R10A),
				.b4(W2R11A),
				.b5(W2R12A),
				.b6(W2R20A),
				.b7(W2R21A),
				.b8(W2R22A),
				.c(c2A01R)
);

ninexnine_unit ninexnine_unit_6879(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2R00B),
				.b1(W2R01B),
				.b2(W2R02B),
				.b3(W2R10B),
				.b4(W2R11B),
				.b5(W2R12B),
				.b6(W2R20B),
				.b7(W2R21B),
				.b8(W2R22B),
				.c(c2B01R)
);

ninexnine_unit ninexnine_unit_6880(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2R00C),
				.b1(W2R01C),
				.b2(W2R02C),
				.b3(W2R10C),
				.b4(W2R11C),
				.b5(W2R12C),
				.b6(W2R20C),
				.b7(W2R21C),
				.b8(W2R22C),
				.c(c2C01R)
);

ninexnine_unit ninexnine_unit_6881(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2R00D),
				.b1(W2R01D),
				.b2(W2R02D),
				.b3(W2R10D),
				.b4(W2R11D),
				.b5(W2R12D),
				.b6(W2R20D),
				.b7(W2R21D),
				.b8(W2R22D),
				.c(c2D01R)
);

ninexnine_unit ninexnine_unit_6882(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2R00E),
				.b1(W2R01E),
				.b2(W2R02E),
				.b3(W2R10E),
				.b4(W2R11E),
				.b5(W2R12E),
				.b6(W2R20E),
				.b7(W2R21E),
				.b8(W2R22E),
				.c(c2E01R)
);

ninexnine_unit ninexnine_unit_6883(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2R00F),
				.b1(W2R01F),
				.b2(W2R02F),
				.b3(W2R10F),
				.b4(W2R11F),
				.b5(W2R12F),
				.b6(W2R20F),
				.b7(W2R21F),
				.b8(W2R22F),
				.c(c2F01R)
);

assign C201R=c2001R+c2101R+c2201R+c2301R+c2401R+c2501R+c2601R+c2701R+c2801R+c2901R+c2A01R+c2B01R+c2C01R+c2D01R+c2E01R+c2F01R;
assign A201R=(C201R>=0)?1:0;

assign P301R=A201R;

ninexnine_unit ninexnine_unit_6884(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2R000),
				.b1(W2R010),
				.b2(W2R020),
				.b3(W2R100),
				.b4(W2R110),
				.b5(W2R120),
				.b6(W2R200),
				.b7(W2R210),
				.b8(W2R220),
				.c(c2002R)
);

ninexnine_unit ninexnine_unit_6885(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2R001),
				.b1(W2R011),
				.b2(W2R021),
				.b3(W2R101),
				.b4(W2R111),
				.b5(W2R121),
				.b6(W2R201),
				.b7(W2R211),
				.b8(W2R221),
				.c(c2102R)
);

ninexnine_unit ninexnine_unit_6886(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2R002),
				.b1(W2R012),
				.b2(W2R022),
				.b3(W2R102),
				.b4(W2R112),
				.b5(W2R122),
				.b6(W2R202),
				.b7(W2R212),
				.b8(W2R222),
				.c(c2202R)
);

ninexnine_unit ninexnine_unit_6887(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2R003),
				.b1(W2R013),
				.b2(W2R023),
				.b3(W2R103),
				.b4(W2R113),
				.b5(W2R123),
				.b6(W2R203),
				.b7(W2R213),
				.b8(W2R223),
				.c(c2302R)
);

ninexnine_unit ninexnine_unit_6888(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2R004),
				.b1(W2R014),
				.b2(W2R024),
				.b3(W2R104),
				.b4(W2R114),
				.b5(W2R124),
				.b6(W2R204),
				.b7(W2R214),
				.b8(W2R224),
				.c(c2402R)
);

ninexnine_unit ninexnine_unit_6889(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2R005),
				.b1(W2R015),
				.b2(W2R025),
				.b3(W2R105),
				.b4(W2R115),
				.b5(W2R125),
				.b6(W2R205),
				.b7(W2R215),
				.b8(W2R225),
				.c(c2502R)
);

ninexnine_unit ninexnine_unit_6890(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2R006),
				.b1(W2R016),
				.b2(W2R026),
				.b3(W2R106),
				.b4(W2R116),
				.b5(W2R126),
				.b6(W2R206),
				.b7(W2R216),
				.b8(W2R226),
				.c(c2602R)
);

ninexnine_unit ninexnine_unit_6891(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2R007),
				.b1(W2R017),
				.b2(W2R027),
				.b3(W2R107),
				.b4(W2R117),
				.b5(W2R127),
				.b6(W2R207),
				.b7(W2R217),
				.b8(W2R227),
				.c(c2702R)
);

ninexnine_unit ninexnine_unit_6892(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2R008),
				.b1(W2R018),
				.b2(W2R028),
				.b3(W2R108),
				.b4(W2R118),
				.b5(W2R128),
				.b6(W2R208),
				.b7(W2R218),
				.b8(W2R228),
				.c(c2802R)
);

ninexnine_unit ninexnine_unit_6893(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2R009),
				.b1(W2R019),
				.b2(W2R029),
				.b3(W2R109),
				.b4(W2R119),
				.b5(W2R129),
				.b6(W2R209),
				.b7(W2R219),
				.b8(W2R229),
				.c(c2902R)
);

ninexnine_unit ninexnine_unit_6894(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2R00A),
				.b1(W2R01A),
				.b2(W2R02A),
				.b3(W2R10A),
				.b4(W2R11A),
				.b5(W2R12A),
				.b6(W2R20A),
				.b7(W2R21A),
				.b8(W2R22A),
				.c(c2A02R)
);

ninexnine_unit ninexnine_unit_6895(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2R00B),
				.b1(W2R01B),
				.b2(W2R02B),
				.b3(W2R10B),
				.b4(W2R11B),
				.b5(W2R12B),
				.b6(W2R20B),
				.b7(W2R21B),
				.b8(W2R22B),
				.c(c2B02R)
);

ninexnine_unit ninexnine_unit_6896(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2R00C),
				.b1(W2R01C),
				.b2(W2R02C),
				.b3(W2R10C),
				.b4(W2R11C),
				.b5(W2R12C),
				.b6(W2R20C),
				.b7(W2R21C),
				.b8(W2R22C),
				.c(c2C02R)
);

ninexnine_unit ninexnine_unit_6897(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2R00D),
				.b1(W2R01D),
				.b2(W2R02D),
				.b3(W2R10D),
				.b4(W2R11D),
				.b5(W2R12D),
				.b6(W2R20D),
				.b7(W2R21D),
				.b8(W2R22D),
				.c(c2D02R)
);

ninexnine_unit ninexnine_unit_6898(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2R00E),
				.b1(W2R01E),
				.b2(W2R02E),
				.b3(W2R10E),
				.b4(W2R11E),
				.b5(W2R12E),
				.b6(W2R20E),
				.b7(W2R21E),
				.b8(W2R22E),
				.c(c2E02R)
);

ninexnine_unit ninexnine_unit_6899(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2R00F),
				.b1(W2R01F),
				.b2(W2R02F),
				.b3(W2R10F),
				.b4(W2R11F),
				.b5(W2R12F),
				.b6(W2R20F),
				.b7(W2R21F),
				.b8(W2R22F),
				.c(c2F02R)
);

assign C202R=c2002R+c2102R+c2202R+c2302R+c2402R+c2502R+c2602R+c2702R+c2802R+c2902R+c2A02R+c2B02R+c2C02R+c2D02R+c2E02R+c2F02R;
assign A202R=(C202R>=0)?1:0;

assign P302R=A202R;

ninexnine_unit ninexnine_unit_6900(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2R000),
				.b1(W2R010),
				.b2(W2R020),
				.b3(W2R100),
				.b4(W2R110),
				.b5(W2R120),
				.b6(W2R200),
				.b7(W2R210),
				.b8(W2R220),
				.c(c2010R)
);

ninexnine_unit ninexnine_unit_6901(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2R001),
				.b1(W2R011),
				.b2(W2R021),
				.b3(W2R101),
				.b4(W2R111),
				.b5(W2R121),
				.b6(W2R201),
				.b7(W2R211),
				.b8(W2R221),
				.c(c2110R)
);

ninexnine_unit ninexnine_unit_6902(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2R002),
				.b1(W2R012),
				.b2(W2R022),
				.b3(W2R102),
				.b4(W2R112),
				.b5(W2R122),
				.b6(W2R202),
				.b7(W2R212),
				.b8(W2R222),
				.c(c2210R)
);

ninexnine_unit ninexnine_unit_6903(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2R003),
				.b1(W2R013),
				.b2(W2R023),
				.b3(W2R103),
				.b4(W2R113),
				.b5(W2R123),
				.b6(W2R203),
				.b7(W2R213),
				.b8(W2R223),
				.c(c2310R)
);

ninexnine_unit ninexnine_unit_6904(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2R004),
				.b1(W2R014),
				.b2(W2R024),
				.b3(W2R104),
				.b4(W2R114),
				.b5(W2R124),
				.b6(W2R204),
				.b7(W2R214),
				.b8(W2R224),
				.c(c2410R)
);

ninexnine_unit ninexnine_unit_6905(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2R005),
				.b1(W2R015),
				.b2(W2R025),
				.b3(W2R105),
				.b4(W2R115),
				.b5(W2R125),
				.b6(W2R205),
				.b7(W2R215),
				.b8(W2R225),
				.c(c2510R)
);

ninexnine_unit ninexnine_unit_6906(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2R006),
				.b1(W2R016),
				.b2(W2R026),
				.b3(W2R106),
				.b4(W2R116),
				.b5(W2R126),
				.b6(W2R206),
				.b7(W2R216),
				.b8(W2R226),
				.c(c2610R)
);

ninexnine_unit ninexnine_unit_6907(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2R007),
				.b1(W2R017),
				.b2(W2R027),
				.b3(W2R107),
				.b4(W2R117),
				.b5(W2R127),
				.b6(W2R207),
				.b7(W2R217),
				.b8(W2R227),
				.c(c2710R)
);

ninexnine_unit ninexnine_unit_6908(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2R008),
				.b1(W2R018),
				.b2(W2R028),
				.b3(W2R108),
				.b4(W2R118),
				.b5(W2R128),
				.b6(W2R208),
				.b7(W2R218),
				.b8(W2R228),
				.c(c2810R)
);

ninexnine_unit ninexnine_unit_6909(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2R009),
				.b1(W2R019),
				.b2(W2R029),
				.b3(W2R109),
				.b4(W2R119),
				.b5(W2R129),
				.b6(W2R209),
				.b7(W2R219),
				.b8(W2R229),
				.c(c2910R)
);

ninexnine_unit ninexnine_unit_6910(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2R00A),
				.b1(W2R01A),
				.b2(W2R02A),
				.b3(W2R10A),
				.b4(W2R11A),
				.b5(W2R12A),
				.b6(W2R20A),
				.b7(W2R21A),
				.b8(W2R22A),
				.c(c2A10R)
);

ninexnine_unit ninexnine_unit_6911(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2R00B),
				.b1(W2R01B),
				.b2(W2R02B),
				.b3(W2R10B),
				.b4(W2R11B),
				.b5(W2R12B),
				.b6(W2R20B),
				.b7(W2R21B),
				.b8(W2R22B),
				.c(c2B10R)
);

ninexnine_unit ninexnine_unit_6912(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2R00C),
				.b1(W2R01C),
				.b2(W2R02C),
				.b3(W2R10C),
				.b4(W2R11C),
				.b5(W2R12C),
				.b6(W2R20C),
				.b7(W2R21C),
				.b8(W2R22C),
				.c(c2C10R)
);

ninexnine_unit ninexnine_unit_6913(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2R00D),
				.b1(W2R01D),
				.b2(W2R02D),
				.b3(W2R10D),
				.b4(W2R11D),
				.b5(W2R12D),
				.b6(W2R20D),
				.b7(W2R21D),
				.b8(W2R22D),
				.c(c2D10R)
);

ninexnine_unit ninexnine_unit_6914(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2R00E),
				.b1(W2R01E),
				.b2(W2R02E),
				.b3(W2R10E),
				.b4(W2R11E),
				.b5(W2R12E),
				.b6(W2R20E),
				.b7(W2R21E),
				.b8(W2R22E),
				.c(c2E10R)
);

ninexnine_unit ninexnine_unit_6915(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2R00F),
				.b1(W2R01F),
				.b2(W2R02F),
				.b3(W2R10F),
				.b4(W2R11F),
				.b5(W2R12F),
				.b6(W2R20F),
				.b7(W2R21F),
				.b8(W2R22F),
				.c(c2F10R)
);

assign C210R=c2010R+c2110R+c2210R+c2310R+c2410R+c2510R+c2610R+c2710R+c2810R+c2910R+c2A10R+c2B10R+c2C10R+c2D10R+c2E10R+c2F10R;
assign A210R=(C210R>=0)?1:0;

assign P310R=A210R;

ninexnine_unit ninexnine_unit_6916(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2R000),
				.b1(W2R010),
				.b2(W2R020),
				.b3(W2R100),
				.b4(W2R110),
				.b5(W2R120),
				.b6(W2R200),
				.b7(W2R210),
				.b8(W2R220),
				.c(c2011R)
);

ninexnine_unit ninexnine_unit_6917(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2R001),
				.b1(W2R011),
				.b2(W2R021),
				.b3(W2R101),
				.b4(W2R111),
				.b5(W2R121),
				.b6(W2R201),
				.b7(W2R211),
				.b8(W2R221),
				.c(c2111R)
);

ninexnine_unit ninexnine_unit_6918(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2R002),
				.b1(W2R012),
				.b2(W2R022),
				.b3(W2R102),
				.b4(W2R112),
				.b5(W2R122),
				.b6(W2R202),
				.b7(W2R212),
				.b8(W2R222),
				.c(c2211R)
);

ninexnine_unit ninexnine_unit_6919(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2R003),
				.b1(W2R013),
				.b2(W2R023),
				.b3(W2R103),
				.b4(W2R113),
				.b5(W2R123),
				.b6(W2R203),
				.b7(W2R213),
				.b8(W2R223),
				.c(c2311R)
);

ninexnine_unit ninexnine_unit_6920(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2R004),
				.b1(W2R014),
				.b2(W2R024),
				.b3(W2R104),
				.b4(W2R114),
				.b5(W2R124),
				.b6(W2R204),
				.b7(W2R214),
				.b8(W2R224),
				.c(c2411R)
);

ninexnine_unit ninexnine_unit_6921(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2R005),
				.b1(W2R015),
				.b2(W2R025),
				.b3(W2R105),
				.b4(W2R115),
				.b5(W2R125),
				.b6(W2R205),
				.b7(W2R215),
				.b8(W2R225),
				.c(c2511R)
);

ninexnine_unit ninexnine_unit_6922(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2R006),
				.b1(W2R016),
				.b2(W2R026),
				.b3(W2R106),
				.b4(W2R116),
				.b5(W2R126),
				.b6(W2R206),
				.b7(W2R216),
				.b8(W2R226),
				.c(c2611R)
);

ninexnine_unit ninexnine_unit_6923(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2R007),
				.b1(W2R017),
				.b2(W2R027),
				.b3(W2R107),
				.b4(W2R117),
				.b5(W2R127),
				.b6(W2R207),
				.b7(W2R217),
				.b8(W2R227),
				.c(c2711R)
);

ninexnine_unit ninexnine_unit_6924(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2R008),
				.b1(W2R018),
				.b2(W2R028),
				.b3(W2R108),
				.b4(W2R118),
				.b5(W2R128),
				.b6(W2R208),
				.b7(W2R218),
				.b8(W2R228),
				.c(c2811R)
);

ninexnine_unit ninexnine_unit_6925(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2R009),
				.b1(W2R019),
				.b2(W2R029),
				.b3(W2R109),
				.b4(W2R119),
				.b5(W2R129),
				.b6(W2R209),
				.b7(W2R219),
				.b8(W2R229),
				.c(c2911R)
);

ninexnine_unit ninexnine_unit_6926(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2R00A),
				.b1(W2R01A),
				.b2(W2R02A),
				.b3(W2R10A),
				.b4(W2R11A),
				.b5(W2R12A),
				.b6(W2R20A),
				.b7(W2R21A),
				.b8(W2R22A),
				.c(c2A11R)
);

ninexnine_unit ninexnine_unit_6927(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2R00B),
				.b1(W2R01B),
				.b2(W2R02B),
				.b3(W2R10B),
				.b4(W2R11B),
				.b5(W2R12B),
				.b6(W2R20B),
				.b7(W2R21B),
				.b8(W2R22B),
				.c(c2B11R)
);

ninexnine_unit ninexnine_unit_6928(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2R00C),
				.b1(W2R01C),
				.b2(W2R02C),
				.b3(W2R10C),
				.b4(W2R11C),
				.b5(W2R12C),
				.b6(W2R20C),
				.b7(W2R21C),
				.b8(W2R22C),
				.c(c2C11R)
);

ninexnine_unit ninexnine_unit_6929(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2R00D),
				.b1(W2R01D),
				.b2(W2R02D),
				.b3(W2R10D),
				.b4(W2R11D),
				.b5(W2R12D),
				.b6(W2R20D),
				.b7(W2R21D),
				.b8(W2R22D),
				.c(c2D11R)
);

ninexnine_unit ninexnine_unit_6930(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2R00E),
				.b1(W2R01E),
				.b2(W2R02E),
				.b3(W2R10E),
				.b4(W2R11E),
				.b5(W2R12E),
				.b6(W2R20E),
				.b7(W2R21E),
				.b8(W2R22E),
				.c(c2E11R)
);

ninexnine_unit ninexnine_unit_6931(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2R00F),
				.b1(W2R01F),
				.b2(W2R02F),
				.b3(W2R10F),
				.b4(W2R11F),
				.b5(W2R12F),
				.b6(W2R20F),
				.b7(W2R21F),
				.b8(W2R22F),
				.c(c2F11R)
);

assign C211R=c2011R+c2111R+c2211R+c2311R+c2411R+c2511R+c2611R+c2711R+c2811R+c2911R+c2A11R+c2B11R+c2C11R+c2D11R+c2E11R+c2F11R;
assign A211R=(C211R>=0)?1:0;

assign P311R=A211R;

ninexnine_unit ninexnine_unit_6932(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2R000),
				.b1(W2R010),
				.b2(W2R020),
				.b3(W2R100),
				.b4(W2R110),
				.b5(W2R120),
				.b6(W2R200),
				.b7(W2R210),
				.b8(W2R220),
				.c(c2012R)
);

ninexnine_unit ninexnine_unit_6933(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2R001),
				.b1(W2R011),
				.b2(W2R021),
				.b3(W2R101),
				.b4(W2R111),
				.b5(W2R121),
				.b6(W2R201),
				.b7(W2R211),
				.b8(W2R221),
				.c(c2112R)
);

ninexnine_unit ninexnine_unit_6934(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2R002),
				.b1(W2R012),
				.b2(W2R022),
				.b3(W2R102),
				.b4(W2R112),
				.b5(W2R122),
				.b6(W2R202),
				.b7(W2R212),
				.b8(W2R222),
				.c(c2212R)
);

ninexnine_unit ninexnine_unit_6935(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2R003),
				.b1(W2R013),
				.b2(W2R023),
				.b3(W2R103),
				.b4(W2R113),
				.b5(W2R123),
				.b6(W2R203),
				.b7(W2R213),
				.b8(W2R223),
				.c(c2312R)
);

ninexnine_unit ninexnine_unit_6936(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2R004),
				.b1(W2R014),
				.b2(W2R024),
				.b3(W2R104),
				.b4(W2R114),
				.b5(W2R124),
				.b6(W2R204),
				.b7(W2R214),
				.b8(W2R224),
				.c(c2412R)
);

ninexnine_unit ninexnine_unit_6937(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2R005),
				.b1(W2R015),
				.b2(W2R025),
				.b3(W2R105),
				.b4(W2R115),
				.b5(W2R125),
				.b6(W2R205),
				.b7(W2R215),
				.b8(W2R225),
				.c(c2512R)
);

ninexnine_unit ninexnine_unit_6938(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2R006),
				.b1(W2R016),
				.b2(W2R026),
				.b3(W2R106),
				.b4(W2R116),
				.b5(W2R126),
				.b6(W2R206),
				.b7(W2R216),
				.b8(W2R226),
				.c(c2612R)
);

ninexnine_unit ninexnine_unit_6939(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2R007),
				.b1(W2R017),
				.b2(W2R027),
				.b3(W2R107),
				.b4(W2R117),
				.b5(W2R127),
				.b6(W2R207),
				.b7(W2R217),
				.b8(W2R227),
				.c(c2712R)
);

ninexnine_unit ninexnine_unit_6940(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2R008),
				.b1(W2R018),
				.b2(W2R028),
				.b3(W2R108),
				.b4(W2R118),
				.b5(W2R128),
				.b6(W2R208),
				.b7(W2R218),
				.b8(W2R228),
				.c(c2812R)
);

ninexnine_unit ninexnine_unit_6941(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2R009),
				.b1(W2R019),
				.b2(W2R029),
				.b3(W2R109),
				.b4(W2R119),
				.b5(W2R129),
				.b6(W2R209),
				.b7(W2R219),
				.b8(W2R229),
				.c(c2912R)
);

ninexnine_unit ninexnine_unit_6942(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2R00A),
				.b1(W2R01A),
				.b2(W2R02A),
				.b3(W2R10A),
				.b4(W2R11A),
				.b5(W2R12A),
				.b6(W2R20A),
				.b7(W2R21A),
				.b8(W2R22A),
				.c(c2A12R)
);

ninexnine_unit ninexnine_unit_6943(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2R00B),
				.b1(W2R01B),
				.b2(W2R02B),
				.b3(W2R10B),
				.b4(W2R11B),
				.b5(W2R12B),
				.b6(W2R20B),
				.b7(W2R21B),
				.b8(W2R22B),
				.c(c2B12R)
);

ninexnine_unit ninexnine_unit_6944(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2R00C),
				.b1(W2R01C),
				.b2(W2R02C),
				.b3(W2R10C),
				.b4(W2R11C),
				.b5(W2R12C),
				.b6(W2R20C),
				.b7(W2R21C),
				.b8(W2R22C),
				.c(c2C12R)
);

ninexnine_unit ninexnine_unit_6945(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2R00D),
				.b1(W2R01D),
				.b2(W2R02D),
				.b3(W2R10D),
				.b4(W2R11D),
				.b5(W2R12D),
				.b6(W2R20D),
				.b7(W2R21D),
				.b8(W2R22D),
				.c(c2D12R)
);

ninexnine_unit ninexnine_unit_6946(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2R00E),
				.b1(W2R01E),
				.b2(W2R02E),
				.b3(W2R10E),
				.b4(W2R11E),
				.b5(W2R12E),
				.b6(W2R20E),
				.b7(W2R21E),
				.b8(W2R22E),
				.c(c2E12R)
);

ninexnine_unit ninexnine_unit_6947(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2R00F),
				.b1(W2R01F),
				.b2(W2R02F),
				.b3(W2R10F),
				.b4(W2R11F),
				.b5(W2R12F),
				.b6(W2R20F),
				.b7(W2R21F),
				.b8(W2R22F),
				.c(c2F12R)
);

assign C212R=c2012R+c2112R+c2212R+c2312R+c2412R+c2512R+c2612R+c2712R+c2812R+c2912R+c2A12R+c2B12R+c2C12R+c2D12R+c2E12R+c2F12R;
assign A212R=(C212R>=0)?1:0;

assign P312R=A212R;

ninexnine_unit ninexnine_unit_6948(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2R000),
				.b1(W2R010),
				.b2(W2R020),
				.b3(W2R100),
				.b4(W2R110),
				.b5(W2R120),
				.b6(W2R200),
				.b7(W2R210),
				.b8(W2R220),
				.c(c2020R)
);

ninexnine_unit ninexnine_unit_6949(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2R001),
				.b1(W2R011),
				.b2(W2R021),
				.b3(W2R101),
				.b4(W2R111),
				.b5(W2R121),
				.b6(W2R201),
				.b7(W2R211),
				.b8(W2R221),
				.c(c2120R)
);

ninexnine_unit ninexnine_unit_6950(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2R002),
				.b1(W2R012),
				.b2(W2R022),
				.b3(W2R102),
				.b4(W2R112),
				.b5(W2R122),
				.b6(W2R202),
				.b7(W2R212),
				.b8(W2R222),
				.c(c2220R)
);

ninexnine_unit ninexnine_unit_6951(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2R003),
				.b1(W2R013),
				.b2(W2R023),
				.b3(W2R103),
				.b4(W2R113),
				.b5(W2R123),
				.b6(W2R203),
				.b7(W2R213),
				.b8(W2R223),
				.c(c2320R)
);

ninexnine_unit ninexnine_unit_6952(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2R004),
				.b1(W2R014),
				.b2(W2R024),
				.b3(W2R104),
				.b4(W2R114),
				.b5(W2R124),
				.b6(W2R204),
				.b7(W2R214),
				.b8(W2R224),
				.c(c2420R)
);

ninexnine_unit ninexnine_unit_6953(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2R005),
				.b1(W2R015),
				.b2(W2R025),
				.b3(W2R105),
				.b4(W2R115),
				.b5(W2R125),
				.b6(W2R205),
				.b7(W2R215),
				.b8(W2R225),
				.c(c2520R)
);

ninexnine_unit ninexnine_unit_6954(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2R006),
				.b1(W2R016),
				.b2(W2R026),
				.b3(W2R106),
				.b4(W2R116),
				.b5(W2R126),
				.b6(W2R206),
				.b7(W2R216),
				.b8(W2R226),
				.c(c2620R)
);

ninexnine_unit ninexnine_unit_6955(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2R007),
				.b1(W2R017),
				.b2(W2R027),
				.b3(W2R107),
				.b4(W2R117),
				.b5(W2R127),
				.b6(W2R207),
				.b7(W2R217),
				.b8(W2R227),
				.c(c2720R)
);

ninexnine_unit ninexnine_unit_6956(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2R008),
				.b1(W2R018),
				.b2(W2R028),
				.b3(W2R108),
				.b4(W2R118),
				.b5(W2R128),
				.b6(W2R208),
				.b7(W2R218),
				.b8(W2R228),
				.c(c2820R)
);

ninexnine_unit ninexnine_unit_6957(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2R009),
				.b1(W2R019),
				.b2(W2R029),
				.b3(W2R109),
				.b4(W2R119),
				.b5(W2R129),
				.b6(W2R209),
				.b7(W2R219),
				.b8(W2R229),
				.c(c2920R)
);

ninexnine_unit ninexnine_unit_6958(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2R00A),
				.b1(W2R01A),
				.b2(W2R02A),
				.b3(W2R10A),
				.b4(W2R11A),
				.b5(W2R12A),
				.b6(W2R20A),
				.b7(W2R21A),
				.b8(W2R22A),
				.c(c2A20R)
);

ninexnine_unit ninexnine_unit_6959(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2R00B),
				.b1(W2R01B),
				.b2(W2R02B),
				.b3(W2R10B),
				.b4(W2R11B),
				.b5(W2R12B),
				.b6(W2R20B),
				.b7(W2R21B),
				.b8(W2R22B),
				.c(c2B20R)
);

ninexnine_unit ninexnine_unit_6960(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2R00C),
				.b1(W2R01C),
				.b2(W2R02C),
				.b3(W2R10C),
				.b4(W2R11C),
				.b5(W2R12C),
				.b6(W2R20C),
				.b7(W2R21C),
				.b8(W2R22C),
				.c(c2C20R)
);

ninexnine_unit ninexnine_unit_6961(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2R00D),
				.b1(W2R01D),
				.b2(W2R02D),
				.b3(W2R10D),
				.b4(W2R11D),
				.b5(W2R12D),
				.b6(W2R20D),
				.b7(W2R21D),
				.b8(W2R22D),
				.c(c2D20R)
);

ninexnine_unit ninexnine_unit_6962(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2R00E),
				.b1(W2R01E),
				.b2(W2R02E),
				.b3(W2R10E),
				.b4(W2R11E),
				.b5(W2R12E),
				.b6(W2R20E),
				.b7(W2R21E),
				.b8(W2R22E),
				.c(c2E20R)
);

ninexnine_unit ninexnine_unit_6963(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2R00F),
				.b1(W2R01F),
				.b2(W2R02F),
				.b3(W2R10F),
				.b4(W2R11F),
				.b5(W2R12F),
				.b6(W2R20F),
				.b7(W2R21F),
				.b8(W2R22F),
				.c(c2F20R)
);

assign C220R=c2020R+c2120R+c2220R+c2320R+c2420R+c2520R+c2620R+c2720R+c2820R+c2920R+c2A20R+c2B20R+c2C20R+c2D20R+c2E20R+c2F20R;
assign A220R=(C220R>=0)?1:0;

assign P320R=A220R;

ninexnine_unit ninexnine_unit_6964(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2R000),
				.b1(W2R010),
				.b2(W2R020),
				.b3(W2R100),
				.b4(W2R110),
				.b5(W2R120),
				.b6(W2R200),
				.b7(W2R210),
				.b8(W2R220),
				.c(c2021R)
);

ninexnine_unit ninexnine_unit_6965(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2R001),
				.b1(W2R011),
				.b2(W2R021),
				.b3(W2R101),
				.b4(W2R111),
				.b5(W2R121),
				.b6(W2R201),
				.b7(W2R211),
				.b8(W2R221),
				.c(c2121R)
);

ninexnine_unit ninexnine_unit_6966(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2R002),
				.b1(W2R012),
				.b2(W2R022),
				.b3(W2R102),
				.b4(W2R112),
				.b5(W2R122),
				.b6(W2R202),
				.b7(W2R212),
				.b8(W2R222),
				.c(c2221R)
);

ninexnine_unit ninexnine_unit_6967(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2R003),
				.b1(W2R013),
				.b2(W2R023),
				.b3(W2R103),
				.b4(W2R113),
				.b5(W2R123),
				.b6(W2R203),
				.b7(W2R213),
				.b8(W2R223),
				.c(c2321R)
);

ninexnine_unit ninexnine_unit_6968(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2R004),
				.b1(W2R014),
				.b2(W2R024),
				.b3(W2R104),
				.b4(W2R114),
				.b5(W2R124),
				.b6(W2R204),
				.b7(W2R214),
				.b8(W2R224),
				.c(c2421R)
);

ninexnine_unit ninexnine_unit_6969(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2R005),
				.b1(W2R015),
				.b2(W2R025),
				.b3(W2R105),
				.b4(W2R115),
				.b5(W2R125),
				.b6(W2R205),
				.b7(W2R215),
				.b8(W2R225),
				.c(c2521R)
);

ninexnine_unit ninexnine_unit_6970(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2R006),
				.b1(W2R016),
				.b2(W2R026),
				.b3(W2R106),
				.b4(W2R116),
				.b5(W2R126),
				.b6(W2R206),
				.b7(W2R216),
				.b8(W2R226),
				.c(c2621R)
);

ninexnine_unit ninexnine_unit_6971(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2R007),
				.b1(W2R017),
				.b2(W2R027),
				.b3(W2R107),
				.b4(W2R117),
				.b5(W2R127),
				.b6(W2R207),
				.b7(W2R217),
				.b8(W2R227),
				.c(c2721R)
);

ninexnine_unit ninexnine_unit_6972(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2R008),
				.b1(W2R018),
				.b2(W2R028),
				.b3(W2R108),
				.b4(W2R118),
				.b5(W2R128),
				.b6(W2R208),
				.b7(W2R218),
				.b8(W2R228),
				.c(c2821R)
);

ninexnine_unit ninexnine_unit_6973(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2R009),
				.b1(W2R019),
				.b2(W2R029),
				.b3(W2R109),
				.b4(W2R119),
				.b5(W2R129),
				.b6(W2R209),
				.b7(W2R219),
				.b8(W2R229),
				.c(c2921R)
);

ninexnine_unit ninexnine_unit_6974(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2R00A),
				.b1(W2R01A),
				.b2(W2R02A),
				.b3(W2R10A),
				.b4(W2R11A),
				.b5(W2R12A),
				.b6(W2R20A),
				.b7(W2R21A),
				.b8(W2R22A),
				.c(c2A21R)
);

ninexnine_unit ninexnine_unit_6975(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2R00B),
				.b1(W2R01B),
				.b2(W2R02B),
				.b3(W2R10B),
				.b4(W2R11B),
				.b5(W2R12B),
				.b6(W2R20B),
				.b7(W2R21B),
				.b8(W2R22B),
				.c(c2B21R)
);

ninexnine_unit ninexnine_unit_6976(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2R00C),
				.b1(W2R01C),
				.b2(W2R02C),
				.b3(W2R10C),
				.b4(W2R11C),
				.b5(W2R12C),
				.b6(W2R20C),
				.b7(W2R21C),
				.b8(W2R22C),
				.c(c2C21R)
);

ninexnine_unit ninexnine_unit_6977(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2R00D),
				.b1(W2R01D),
				.b2(W2R02D),
				.b3(W2R10D),
				.b4(W2R11D),
				.b5(W2R12D),
				.b6(W2R20D),
				.b7(W2R21D),
				.b8(W2R22D),
				.c(c2D21R)
);

ninexnine_unit ninexnine_unit_6978(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2R00E),
				.b1(W2R01E),
				.b2(W2R02E),
				.b3(W2R10E),
				.b4(W2R11E),
				.b5(W2R12E),
				.b6(W2R20E),
				.b7(W2R21E),
				.b8(W2R22E),
				.c(c2E21R)
);

ninexnine_unit ninexnine_unit_6979(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2R00F),
				.b1(W2R01F),
				.b2(W2R02F),
				.b3(W2R10F),
				.b4(W2R11F),
				.b5(W2R12F),
				.b6(W2R20F),
				.b7(W2R21F),
				.b8(W2R22F),
				.c(c2F21R)
);

assign C221R=c2021R+c2121R+c2221R+c2321R+c2421R+c2521R+c2621R+c2721R+c2821R+c2921R+c2A21R+c2B21R+c2C21R+c2D21R+c2E21R+c2F21R;
assign A221R=(C221R>=0)?1:0;

assign P321R=A221R;

ninexnine_unit ninexnine_unit_6980(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2R000),
				.b1(W2R010),
				.b2(W2R020),
				.b3(W2R100),
				.b4(W2R110),
				.b5(W2R120),
				.b6(W2R200),
				.b7(W2R210),
				.b8(W2R220),
				.c(c2022R)
);

ninexnine_unit ninexnine_unit_6981(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2R001),
				.b1(W2R011),
				.b2(W2R021),
				.b3(W2R101),
				.b4(W2R111),
				.b5(W2R121),
				.b6(W2R201),
				.b7(W2R211),
				.b8(W2R221),
				.c(c2122R)
);

ninexnine_unit ninexnine_unit_6982(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2R002),
				.b1(W2R012),
				.b2(W2R022),
				.b3(W2R102),
				.b4(W2R112),
				.b5(W2R122),
				.b6(W2R202),
				.b7(W2R212),
				.b8(W2R222),
				.c(c2222R)
);

ninexnine_unit ninexnine_unit_6983(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2R003),
				.b1(W2R013),
				.b2(W2R023),
				.b3(W2R103),
				.b4(W2R113),
				.b5(W2R123),
				.b6(W2R203),
				.b7(W2R213),
				.b8(W2R223),
				.c(c2322R)
);

ninexnine_unit ninexnine_unit_6984(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2R004),
				.b1(W2R014),
				.b2(W2R024),
				.b3(W2R104),
				.b4(W2R114),
				.b5(W2R124),
				.b6(W2R204),
				.b7(W2R214),
				.b8(W2R224),
				.c(c2422R)
);

ninexnine_unit ninexnine_unit_6985(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2R005),
				.b1(W2R015),
				.b2(W2R025),
				.b3(W2R105),
				.b4(W2R115),
				.b5(W2R125),
				.b6(W2R205),
				.b7(W2R215),
				.b8(W2R225),
				.c(c2522R)
);

ninexnine_unit ninexnine_unit_6986(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2R006),
				.b1(W2R016),
				.b2(W2R026),
				.b3(W2R106),
				.b4(W2R116),
				.b5(W2R126),
				.b6(W2R206),
				.b7(W2R216),
				.b8(W2R226),
				.c(c2622R)
);

ninexnine_unit ninexnine_unit_6987(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2R007),
				.b1(W2R017),
				.b2(W2R027),
				.b3(W2R107),
				.b4(W2R117),
				.b5(W2R127),
				.b6(W2R207),
				.b7(W2R217),
				.b8(W2R227),
				.c(c2722R)
);

ninexnine_unit ninexnine_unit_6988(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2R008),
				.b1(W2R018),
				.b2(W2R028),
				.b3(W2R108),
				.b4(W2R118),
				.b5(W2R128),
				.b6(W2R208),
				.b7(W2R218),
				.b8(W2R228),
				.c(c2822R)
);

ninexnine_unit ninexnine_unit_6989(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2R009),
				.b1(W2R019),
				.b2(W2R029),
				.b3(W2R109),
				.b4(W2R119),
				.b5(W2R129),
				.b6(W2R209),
				.b7(W2R219),
				.b8(W2R229),
				.c(c2922R)
);

ninexnine_unit ninexnine_unit_6990(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2R00A),
				.b1(W2R01A),
				.b2(W2R02A),
				.b3(W2R10A),
				.b4(W2R11A),
				.b5(W2R12A),
				.b6(W2R20A),
				.b7(W2R21A),
				.b8(W2R22A),
				.c(c2A22R)
);

ninexnine_unit ninexnine_unit_6991(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2R00B),
				.b1(W2R01B),
				.b2(W2R02B),
				.b3(W2R10B),
				.b4(W2R11B),
				.b5(W2R12B),
				.b6(W2R20B),
				.b7(W2R21B),
				.b8(W2R22B),
				.c(c2B22R)
);

ninexnine_unit ninexnine_unit_6992(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2R00C),
				.b1(W2R01C),
				.b2(W2R02C),
				.b3(W2R10C),
				.b4(W2R11C),
				.b5(W2R12C),
				.b6(W2R20C),
				.b7(W2R21C),
				.b8(W2R22C),
				.c(c2C22R)
);

ninexnine_unit ninexnine_unit_6993(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2R00D),
				.b1(W2R01D),
				.b2(W2R02D),
				.b3(W2R10D),
				.b4(W2R11D),
				.b5(W2R12D),
				.b6(W2R20D),
				.b7(W2R21D),
				.b8(W2R22D),
				.c(c2D22R)
);

ninexnine_unit ninexnine_unit_6994(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2R00E),
				.b1(W2R01E),
				.b2(W2R02E),
				.b3(W2R10E),
				.b4(W2R11E),
				.b5(W2R12E),
				.b6(W2R20E),
				.b7(W2R21E),
				.b8(W2R22E),
				.c(c2E22R)
);

ninexnine_unit ninexnine_unit_6995(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2R00F),
				.b1(W2R01F),
				.b2(W2R02F),
				.b3(W2R10F),
				.b4(W2R11F),
				.b5(W2R12F),
				.b6(W2R20F),
				.b7(W2R21F),
				.b8(W2R22F),
				.c(c2F22R)
);

assign C222R=c2022R+c2122R+c2222R+c2322R+c2422R+c2522R+c2622R+c2722R+c2822R+c2922R+c2A22R+c2B22R+c2C22R+c2D22R+c2E22R+c2F22R;
assign A222R=(C222R>=0)?1:0;

assign P322R=A222R;

ninexnine_unit ninexnine_unit_6996(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2S000),
				.b1(W2S010),
				.b2(W2S020),
				.b3(W2S100),
				.b4(W2S110),
				.b5(W2S120),
				.b6(W2S200),
				.b7(W2S210),
				.b8(W2S220),
				.c(c2000S)
);

ninexnine_unit ninexnine_unit_6997(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2S001),
				.b1(W2S011),
				.b2(W2S021),
				.b3(W2S101),
				.b4(W2S111),
				.b5(W2S121),
				.b6(W2S201),
				.b7(W2S211),
				.b8(W2S221),
				.c(c2100S)
);

ninexnine_unit ninexnine_unit_6998(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2S002),
				.b1(W2S012),
				.b2(W2S022),
				.b3(W2S102),
				.b4(W2S112),
				.b5(W2S122),
				.b6(W2S202),
				.b7(W2S212),
				.b8(W2S222),
				.c(c2200S)
);

ninexnine_unit ninexnine_unit_6999(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2S003),
				.b1(W2S013),
				.b2(W2S023),
				.b3(W2S103),
				.b4(W2S113),
				.b5(W2S123),
				.b6(W2S203),
				.b7(W2S213),
				.b8(W2S223),
				.c(c2300S)
);

ninexnine_unit ninexnine_unit_7000(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2S004),
				.b1(W2S014),
				.b2(W2S024),
				.b3(W2S104),
				.b4(W2S114),
				.b5(W2S124),
				.b6(W2S204),
				.b7(W2S214),
				.b8(W2S224),
				.c(c2400S)
);

ninexnine_unit ninexnine_unit_7001(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2S005),
				.b1(W2S015),
				.b2(W2S025),
				.b3(W2S105),
				.b4(W2S115),
				.b5(W2S125),
				.b6(W2S205),
				.b7(W2S215),
				.b8(W2S225),
				.c(c2500S)
);

ninexnine_unit ninexnine_unit_7002(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2S006),
				.b1(W2S016),
				.b2(W2S026),
				.b3(W2S106),
				.b4(W2S116),
				.b5(W2S126),
				.b6(W2S206),
				.b7(W2S216),
				.b8(W2S226),
				.c(c2600S)
);

ninexnine_unit ninexnine_unit_7003(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2S007),
				.b1(W2S017),
				.b2(W2S027),
				.b3(W2S107),
				.b4(W2S117),
				.b5(W2S127),
				.b6(W2S207),
				.b7(W2S217),
				.b8(W2S227),
				.c(c2700S)
);

ninexnine_unit ninexnine_unit_7004(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2S008),
				.b1(W2S018),
				.b2(W2S028),
				.b3(W2S108),
				.b4(W2S118),
				.b5(W2S128),
				.b6(W2S208),
				.b7(W2S218),
				.b8(W2S228),
				.c(c2800S)
);

ninexnine_unit ninexnine_unit_7005(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2S009),
				.b1(W2S019),
				.b2(W2S029),
				.b3(W2S109),
				.b4(W2S119),
				.b5(W2S129),
				.b6(W2S209),
				.b7(W2S219),
				.b8(W2S229),
				.c(c2900S)
);

ninexnine_unit ninexnine_unit_7006(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2S00A),
				.b1(W2S01A),
				.b2(W2S02A),
				.b3(W2S10A),
				.b4(W2S11A),
				.b5(W2S12A),
				.b6(W2S20A),
				.b7(W2S21A),
				.b8(W2S22A),
				.c(c2A00S)
);

ninexnine_unit ninexnine_unit_7007(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2S00B),
				.b1(W2S01B),
				.b2(W2S02B),
				.b3(W2S10B),
				.b4(W2S11B),
				.b5(W2S12B),
				.b6(W2S20B),
				.b7(W2S21B),
				.b8(W2S22B),
				.c(c2B00S)
);

ninexnine_unit ninexnine_unit_7008(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2S00C),
				.b1(W2S01C),
				.b2(W2S02C),
				.b3(W2S10C),
				.b4(W2S11C),
				.b5(W2S12C),
				.b6(W2S20C),
				.b7(W2S21C),
				.b8(W2S22C),
				.c(c2C00S)
);

ninexnine_unit ninexnine_unit_7009(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2S00D),
				.b1(W2S01D),
				.b2(W2S02D),
				.b3(W2S10D),
				.b4(W2S11D),
				.b5(W2S12D),
				.b6(W2S20D),
				.b7(W2S21D),
				.b8(W2S22D),
				.c(c2D00S)
);

ninexnine_unit ninexnine_unit_7010(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2S00E),
				.b1(W2S01E),
				.b2(W2S02E),
				.b3(W2S10E),
				.b4(W2S11E),
				.b5(W2S12E),
				.b6(W2S20E),
				.b7(W2S21E),
				.b8(W2S22E),
				.c(c2E00S)
);

ninexnine_unit ninexnine_unit_7011(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2S00F),
				.b1(W2S01F),
				.b2(W2S02F),
				.b3(W2S10F),
				.b4(W2S11F),
				.b5(W2S12F),
				.b6(W2S20F),
				.b7(W2S21F),
				.b8(W2S22F),
				.c(c2F00S)
);

assign C200S=c2000S+c2100S+c2200S+c2300S+c2400S+c2500S+c2600S+c2700S+c2800S+c2900S+c2A00S+c2B00S+c2C00S+c2D00S+c2E00S+c2F00S;
assign A200S=(C200S>=0)?1:0;

assign P300S=A200S;

ninexnine_unit ninexnine_unit_7012(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2S000),
				.b1(W2S010),
				.b2(W2S020),
				.b3(W2S100),
				.b4(W2S110),
				.b5(W2S120),
				.b6(W2S200),
				.b7(W2S210),
				.b8(W2S220),
				.c(c2001S)
);

ninexnine_unit ninexnine_unit_7013(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2S001),
				.b1(W2S011),
				.b2(W2S021),
				.b3(W2S101),
				.b4(W2S111),
				.b5(W2S121),
				.b6(W2S201),
				.b7(W2S211),
				.b8(W2S221),
				.c(c2101S)
);

ninexnine_unit ninexnine_unit_7014(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2S002),
				.b1(W2S012),
				.b2(W2S022),
				.b3(W2S102),
				.b4(W2S112),
				.b5(W2S122),
				.b6(W2S202),
				.b7(W2S212),
				.b8(W2S222),
				.c(c2201S)
);

ninexnine_unit ninexnine_unit_7015(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2S003),
				.b1(W2S013),
				.b2(W2S023),
				.b3(W2S103),
				.b4(W2S113),
				.b5(W2S123),
				.b6(W2S203),
				.b7(W2S213),
				.b8(W2S223),
				.c(c2301S)
);

ninexnine_unit ninexnine_unit_7016(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2S004),
				.b1(W2S014),
				.b2(W2S024),
				.b3(W2S104),
				.b4(W2S114),
				.b5(W2S124),
				.b6(W2S204),
				.b7(W2S214),
				.b8(W2S224),
				.c(c2401S)
);

ninexnine_unit ninexnine_unit_7017(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2S005),
				.b1(W2S015),
				.b2(W2S025),
				.b3(W2S105),
				.b4(W2S115),
				.b5(W2S125),
				.b6(W2S205),
				.b7(W2S215),
				.b8(W2S225),
				.c(c2501S)
);

ninexnine_unit ninexnine_unit_7018(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2S006),
				.b1(W2S016),
				.b2(W2S026),
				.b3(W2S106),
				.b4(W2S116),
				.b5(W2S126),
				.b6(W2S206),
				.b7(W2S216),
				.b8(W2S226),
				.c(c2601S)
);

ninexnine_unit ninexnine_unit_7019(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2S007),
				.b1(W2S017),
				.b2(W2S027),
				.b3(W2S107),
				.b4(W2S117),
				.b5(W2S127),
				.b6(W2S207),
				.b7(W2S217),
				.b8(W2S227),
				.c(c2701S)
);

ninexnine_unit ninexnine_unit_7020(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2S008),
				.b1(W2S018),
				.b2(W2S028),
				.b3(W2S108),
				.b4(W2S118),
				.b5(W2S128),
				.b6(W2S208),
				.b7(W2S218),
				.b8(W2S228),
				.c(c2801S)
);

ninexnine_unit ninexnine_unit_7021(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2S009),
				.b1(W2S019),
				.b2(W2S029),
				.b3(W2S109),
				.b4(W2S119),
				.b5(W2S129),
				.b6(W2S209),
				.b7(W2S219),
				.b8(W2S229),
				.c(c2901S)
);

ninexnine_unit ninexnine_unit_7022(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2S00A),
				.b1(W2S01A),
				.b2(W2S02A),
				.b3(W2S10A),
				.b4(W2S11A),
				.b5(W2S12A),
				.b6(W2S20A),
				.b7(W2S21A),
				.b8(W2S22A),
				.c(c2A01S)
);

ninexnine_unit ninexnine_unit_7023(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2S00B),
				.b1(W2S01B),
				.b2(W2S02B),
				.b3(W2S10B),
				.b4(W2S11B),
				.b5(W2S12B),
				.b6(W2S20B),
				.b7(W2S21B),
				.b8(W2S22B),
				.c(c2B01S)
);

ninexnine_unit ninexnine_unit_7024(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2S00C),
				.b1(W2S01C),
				.b2(W2S02C),
				.b3(W2S10C),
				.b4(W2S11C),
				.b5(W2S12C),
				.b6(W2S20C),
				.b7(W2S21C),
				.b8(W2S22C),
				.c(c2C01S)
);

ninexnine_unit ninexnine_unit_7025(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2S00D),
				.b1(W2S01D),
				.b2(W2S02D),
				.b3(W2S10D),
				.b4(W2S11D),
				.b5(W2S12D),
				.b6(W2S20D),
				.b7(W2S21D),
				.b8(W2S22D),
				.c(c2D01S)
);

ninexnine_unit ninexnine_unit_7026(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2S00E),
				.b1(W2S01E),
				.b2(W2S02E),
				.b3(W2S10E),
				.b4(W2S11E),
				.b5(W2S12E),
				.b6(W2S20E),
				.b7(W2S21E),
				.b8(W2S22E),
				.c(c2E01S)
);

ninexnine_unit ninexnine_unit_7027(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2S00F),
				.b1(W2S01F),
				.b2(W2S02F),
				.b3(W2S10F),
				.b4(W2S11F),
				.b5(W2S12F),
				.b6(W2S20F),
				.b7(W2S21F),
				.b8(W2S22F),
				.c(c2F01S)
);

assign C201S=c2001S+c2101S+c2201S+c2301S+c2401S+c2501S+c2601S+c2701S+c2801S+c2901S+c2A01S+c2B01S+c2C01S+c2D01S+c2E01S+c2F01S;
assign A201S=(C201S>=0)?1:0;

assign P301S=A201S;

ninexnine_unit ninexnine_unit_7028(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2S000),
				.b1(W2S010),
				.b2(W2S020),
				.b3(W2S100),
				.b4(W2S110),
				.b5(W2S120),
				.b6(W2S200),
				.b7(W2S210),
				.b8(W2S220),
				.c(c2002S)
);

ninexnine_unit ninexnine_unit_7029(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2S001),
				.b1(W2S011),
				.b2(W2S021),
				.b3(W2S101),
				.b4(W2S111),
				.b5(W2S121),
				.b6(W2S201),
				.b7(W2S211),
				.b8(W2S221),
				.c(c2102S)
);

ninexnine_unit ninexnine_unit_7030(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2S002),
				.b1(W2S012),
				.b2(W2S022),
				.b3(W2S102),
				.b4(W2S112),
				.b5(W2S122),
				.b6(W2S202),
				.b7(W2S212),
				.b8(W2S222),
				.c(c2202S)
);

ninexnine_unit ninexnine_unit_7031(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2S003),
				.b1(W2S013),
				.b2(W2S023),
				.b3(W2S103),
				.b4(W2S113),
				.b5(W2S123),
				.b6(W2S203),
				.b7(W2S213),
				.b8(W2S223),
				.c(c2302S)
);

ninexnine_unit ninexnine_unit_7032(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2S004),
				.b1(W2S014),
				.b2(W2S024),
				.b3(W2S104),
				.b4(W2S114),
				.b5(W2S124),
				.b6(W2S204),
				.b7(W2S214),
				.b8(W2S224),
				.c(c2402S)
);

ninexnine_unit ninexnine_unit_7033(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2S005),
				.b1(W2S015),
				.b2(W2S025),
				.b3(W2S105),
				.b4(W2S115),
				.b5(W2S125),
				.b6(W2S205),
				.b7(W2S215),
				.b8(W2S225),
				.c(c2502S)
);

ninexnine_unit ninexnine_unit_7034(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2S006),
				.b1(W2S016),
				.b2(W2S026),
				.b3(W2S106),
				.b4(W2S116),
				.b5(W2S126),
				.b6(W2S206),
				.b7(W2S216),
				.b8(W2S226),
				.c(c2602S)
);

ninexnine_unit ninexnine_unit_7035(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2S007),
				.b1(W2S017),
				.b2(W2S027),
				.b3(W2S107),
				.b4(W2S117),
				.b5(W2S127),
				.b6(W2S207),
				.b7(W2S217),
				.b8(W2S227),
				.c(c2702S)
);

ninexnine_unit ninexnine_unit_7036(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2S008),
				.b1(W2S018),
				.b2(W2S028),
				.b3(W2S108),
				.b4(W2S118),
				.b5(W2S128),
				.b6(W2S208),
				.b7(W2S218),
				.b8(W2S228),
				.c(c2802S)
);

ninexnine_unit ninexnine_unit_7037(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2S009),
				.b1(W2S019),
				.b2(W2S029),
				.b3(W2S109),
				.b4(W2S119),
				.b5(W2S129),
				.b6(W2S209),
				.b7(W2S219),
				.b8(W2S229),
				.c(c2902S)
);

ninexnine_unit ninexnine_unit_7038(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2S00A),
				.b1(W2S01A),
				.b2(W2S02A),
				.b3(W2S10A),
				.b4(W2S11A),
				.b5(W2S12A),
				.b6(W2S20A),
				.b7(W2S21A),
				.b8(W2S22A),
				.c(c2A02S)
);

ninexnine_unit ninexnine_unit_7039(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2S00B),
				.b1(W2S01B),
				.b2(W2S02B),
				.b3(W2S10B),
				.b4(W2S11B),
				.b5(W2S12B),
				.b6(W2S20B),
				.b7(W2S21B),
				.b8(W2S22B),
				.c(c2B02S)
);

ninexnine_unit ninexnine_unit_7040(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2S00C),
				.b1(W2S01C),
				.b2(W2S02C),
				.b3(W2S10C),
				.b4(W2S11C),
				.b5(W2S12C),
				.b6(W2S20C),
				.b7(W2S21C),
				.b8(W2S22C),
				.c(c2C02S)
);

ninexnine_unit ninexnine_unit_7041(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2S00D),
				.b1(W2S01D),
				.b2(W2S02D),
				.b3(W2S10D),
				.b4(W2S11D),
				.b5(W2S12D),
				.b6(W2S20D),
				.b7(W2S21D),
				.b8(W2S22D),
				.c(c2D02S)
);

ninexnine_unit ninexnine_unit_7042(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2S00E),
				.b1(W2S01E),
				.b2(W2S02E),
				.b3(W2S10E),
				.b4(W2S11E),
				.b5(W2S12E),
				.b6(W2S20E),
				.b7(W2S21E),
				.b8(W2S22E),
				.c(c2E02S)
);

ninexnine_unit ninexnine_unit_7043(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2S00F),
				.b1(W2S01F),
				.b2(W2S02F),
				.b3(W2S10F),
				.b4(W2S11F),
				.b5(W2S12F),
				.b6(W2S20F),
				.b7(W2S21F),
				.b8(W2S22F),
				.c(c2F02S)
);

assign C202S=c2002S+c2102S+c2202S+c2302S+c2402S+c2502S+c2602S+c2702S+c2802S+c2902S+c2A02S+c2B02S+c2C02S+c2D02S+c2E02S+c2F02S;
assign A202S=(C202S>=0)?1:0;

assign P302S=A202S;

ninexnine_unit ninexnine_unit_7044(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2S000),
				.b1(W2S010),
				.b2(W2S020),
				.b3(W2S100),
				.b4(W2S110),
				.b5(W2S120),
				.b6(W2S200),
				.b7(W2S210),
				.b8(W2S220),
				.c(c2010S)
);

ninexnine_unit ninexnine_unit_7045(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2S001),
				.b1(W2S011),
				.b2(W2S021),
				.b3(W2S101),
				.b4(W2S111),
				.b5(W2S121),
				.b6(W2S201),
				.b7(W2S211),
				.b8(W2S221),
				.c(c2110S)
);

ninexnine_unit ninexnine_unit_7046(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2S002),
				.b1(W2S012),
				.b2(W2S022),
				.b3(W2S102),
				.b4(W2S112),
				.b5(W2S122),
				.b6(W2S202),
				.b7(W2S212),
				.b8(W2S222),
				.c(c2210S)
);

ninexnine_unit ninexnine_unit_7047(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2S003),
				.b1(W2S013),
				.b2(W2S023),
				.b3(W2S103),
				.b4(W2S113),
				.b5(W2S123),
				.b6(W2S203),
				.b7(W2S213),
				.b8(W2S223),
				.c(c2310S)
);

ninexnine_unit ninexnine_unit_7048(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2S004),
				.b1(W2S014),
				.b2(W2S024),
				.b3(W2S104),
				.b4(W2S114),
				.b5(W2S124),
				.b6(W2S204),
				.b7(W2S214),
				.b8(W2S224),
				.c(c2410S)
);

ninexnine_unit ninexnine_unit_7049(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2S005),
				.b1(W2S015),
				.b2(W2S025),
				.b3(W2S105),
				.b4(W2S115),
				.b5(W2S125),
				.b6(W2S205),
				.b7(W2S215),
				.b8(W2S225),
				.c(c2510S)
);

ninexnine_unit ninexnine_unit_7050(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2S006),
				.b1(W2S016),
				.b2(W2S026),
				.b3(W2S106),
				.b4(W2S116),
				.b5(W2S126),
				.b6(W2S206),
				.b7(W2S216),
				.b8(W2S226),
				.c(c2610S)
);

ninexnine_unit ninexnine_unit_7051(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2S007),
				.b1(W2S017),
				.b2(W2S027),
				.b3(W2S107),
				.b4(W2S117),
				.b5(W2S127),
				.b6(W2S207),
				.b7(W2S217),
				.b8(W2S227),
				.c(c2710S)
);

ninexnine_unit ninexnine_unit_7052(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2S008),
				.b1(W2S018),
				.b2(W2S028),
				.b3(W2S108),
				.b4(W2S118),
				.b5(W2S128),
				.b6(W2S208),
				.b7(W2S218),
				.b8(W2S228),
				.c(c2810S)
);

ninexnine_unit ninexnine_unit_7053(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2S009),
				.b1(W2S019),
				.b2(W2S029),
				.b3(W2S109),
				.b4(W2S119),
				.b5(W2S129),
				.b6(W2S209),
				.b7(W2S219),
				.b8(W2S229),
				.c(c2910S)
);

ninexnine_unit ninexnine_unit_7054(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2S00A),
				.b1(W2S01A),
				.b2(W2S02A),
				.b3(W2S10A),
				.b4(W2S11A),
				.b5(W2S12A),
				.b6(W2S20A),
				.b7(W2S21A),
				.b8(W2S22A),
				.c(c2A10S)
);

ninexnine_unit ninexnine_unit_7055(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2S00B),
				.b1(W2S01B),
				.b2(W2S02B),
				.b3(W2S10B),
				.b4(W2S11B),
				.b5(W2S12B),
				.b6(W2S20B),
				.b7(W2S21B),
				.b8(W2S22B),
				.c(c2B10S)
);

ninexnine_unit ninexnine_unit_7056(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2S00C),
				.b1(W2S01C),
				.b2(W2S02C),
				.b3(W2S10C),
				.b4(W2S11C),
				.b5(W2S12C),
				.b6(W2S20C),
				.b7(W2S21C),
				.b8(W2S22C),
				.c(c2C10S)
);

ninexnine_unit ninexnine_unit_7057(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2S00D),
				.b1(W2S01D),
				.b2(W2S02D),
				.b3(W2S10D),
				.b4(W2S11D),
				.b5(W2S12D),
				.b6(W2S20D),
				.b7(W2S21D),
				.b8(W2S22D),
				.c(c2D10S)
);

ninexnine_unit ninexnine_unit_7058(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2S00E),
				.b1(W2S01E),
				.b2(W2S02E),
				.b3(W2S10E),
				.b4(W2S11E),
				.b5(W2S12E),
				.b6(W2S20E),
				.b7(W2S21E),
				.b8(W2S22E),
				.c(c2E10S)
);

ninexnine_unit ninexnine_unit_7059(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2S00F),
				.b1(W2S01F),
				.b2(W2S02F),
				.b3(W2S10F),
				.b4(W2S11F),
				.b5(W2S12F),
				.b6(W2S20F),
				.b7(W2S21F),
				.b8(W2S22F),
				.c(c2F10S)
);

assign C210S=c2010S+c2110S+c2210S+c2310S+c2410S+c2510S+c2610S+c2710S+c2810S+c2910S+c2A10S+c2B10S+c2C10S+c2D10S+c2E10S+c2F10S;
assign A210S=(C210S>=0)?1:0;

assign P310S=A210S;

ninexnine_unit ninexnine_unit_7060(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2S000),
				.b1(W2S010),
				.b2(W2S020),
				.b3(W2S100),
				.b4(W2S110),
				.b5(W2S120),
				.b6(W2S200),
				.b7(W2S210),
				.b8(W2S220),
				.c(c2011S)
);

ninexnine_unit ninexnine_unit_7061(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2S001),
				.b1(W2S011),
				.b2(W2S021),
				.b3(W2S101),
				.b4(W2S111),
				.b5(W2S121),
				.b6(W2S201),
				.b7(W2S211),
				.b8(W2S221),
				.c(c2111S)
);

ninexnine_unit ninexnine_unit_7062(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2S002),
				.b1(W2S012),
				.b2(W2S022),
				.b3(W2S102),
				.b4(W2S112),
				.b5(W2S122),
				.b6(W2S202),
				.b7(W2S212),
				.b8(W2S222),
				.c(c2211S)
);

ninexnine_unit ninexnine_unit_7063(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2S003),
				.b1(W2S013),
				.b2(W2S023),
				.b3(W2S103),
				.b4(W2S113),
				.b5(W2S123),
				.b6(W2S203),
				.b7(W2S213),
				.b8(W2S223),
				.c(c2311S)
);

ninexnine_unit ninexnine_unit_7064(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2S004),
				.b1(W2S014),
				.b2(W2S024),
				.b3(W2S104),
				.b4(W2S114),
				.b5(W2S124),
				.b6(W2S204),
				.b7(W2S214),
				.b8(W2S224),
				.c(c2411S)
);

ninexnine_unit ninexnine_unit_7065(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2S005),
				.b1(W2S015),
				.b2(W2S025),
				.b3(W2S105),
				.b4(W2S115),
				.b5(W2S125),
				.b6(W2S205),
				.b7(W2S215),
				.b8(W2S225),
				.c(c2511S)
);

ninexnine_unit ninexnine_unit_7066(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2S006),
				.b1(W2S016),
				.b2(W2S026),
				.b3(W2S106),
				.b4(W2S116),
				.b5(W2S126),
				.b6(W2S206),
				.b7(W2S216),
				.b8(W2S226),
				.c(c2611S)
);

ninexnine_unit ninexnine_unit_7067(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2S007),
				.b1(W2S017),
				.b2(W2S027),
				.b3(W2S107),
				.b4(W2S117),
				.b5(W2S127),
				.b6(W2S207),
				.b7(W2S217),
				.b8(W2S227),
				.c(c2711S)
);

ninexnine_unit ninexnine_unit_7068(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2S008),
				.b1(W2S018),
				.b2(W2S028),
				.b3(W2S108),
				.b4(W2S118),
				.b5(W2S128),
				.b6(W2S208),
				.b7(W2S218),
				.b8(W2S228),
				.c(c2811S)
);

ninexnine_unit ninexnine_unit_7069(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2S009),
				.b1(W2S019),
				.b2(W2S029),
				.b3(W2S109),
				.b4(W2S119),
				.b5(W2S129),
				.b6(W2S209),
				.b7(W2S219),
				.b8(W2S229),
				.c(c2911S)
);

ninexnine_unit ninexnine_unit_7070(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2S00A),
				.b1(W2S01A),
				.b2(W2S02A),
				.b3(W2S10A),
				.b4(W2S11A),
				.b5(W2S12A),
				.b6(W2S20A),
				.b7(W2S21A),
				.b8(W2S22A),
				.c(c2A11S)
);

ninexnine_unit ninexnine_unit_7071(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2S00B),
				.b1(W2S01B),
				.b2(W2S02B),
				.b3(W2S10B),
				.b4(W2S11B),
				.b5(W2S12B),
				.b6(W2S20B),
				.b7(W2S21B),
				.b8(W2S22B),
				.c(c2B11S)
);

ninexnine_unit ninexnine_unit_7072(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2S00C),
				.b1(W2S01C),
				.b2(W2S02C),
				.b3(W2S10C),
				.b4(W2S11C),
				.b5(W2S12C),
				.b6(W2S20C),
				.b7(W2S21C),
				.b8(W2S22C),
				.c(c2C11S)
);

ninexnine_unit ninexnine_unit_7073(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2S00D),
				.b1(W2S01D),
				.b2(W2S02D),
				.b3(W2S10D),
				.b4(W2S11D),
				.b5(W2S12D),
				.b6(W2S20D),
				.b7(W2S21D),
				.b8(W2S22D),
				.c(c2D11S)
);

ninexnine_unit ninexnine_unit_7074(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2S00E),
				.b1(W2S01E),
				.b2(W2S02E),
				.b3(W2S10E),
				.b4(W2S11E),
				.b5(W2S12E),
				.b6(W2S20E),
				.b7(W2S21E),
				.b8(W2S22E),
				.c(c2E11S)
);

ninexnine_unit ninexnine_unit_7075(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2S00F),
				.b1(W2S01F),
				.b2(W2S02F),
				.b3(W2S10F),
				.b4(W2S11F),
				.b5(W2S12F),
				.b6(W2S20F),
				.b7(W2S21F),
				.b8(W2S22F),
				.c(c2F11S)
);

assign C211S=c2011S+c2111S+c2211S+c2311S+c2411S+c2511S+c2611S+c2711S+c2811S+c2911S+c2A11S+c2B11S+c2C11S+c2D11S+c2E11S+c2F11S;
assign A211S=(C211S>=0)?1:0;

assign P311S=A211S;

ninexnine_unit ninexnine_unit_7076(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2S000),
				.b1(W2S010),
				.b2(W2S020),
				.b3(W2S100),
				.b4(W2S110),
				.b5(W2S120),
				.b6(W2S200),
				.b7(W2S210),
				.b8(W2S220),
				.c(c2012S)
);

ninexnine_unit ninexnine_unit_7077(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2S001),
				.b1(W2S011),
				.b2(W2S021),
				.b3(W2S101),
				.b4(W2S111),
				.b5(W2S121),
				.b6(W2S201),
				.b7(W2S211),
				.b8(W2S221),
				.c(c2112S)
);

ninexnine_unit ninexnine_unit_7078(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2S002),
				.b1(W2S012),
				.b2(W2S022),
				.b3(W2S102),
				.b4(W2S112),
				.b5(W2S122),
				.b6(W2S202),
				.b7(W2S212),
				.b8(W2S222),
				.c(c2212S)
);

ninexnine_unit ninexnine_unit_7079(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2S003),
				.b1(W2S013),
				.b2(W2S023),
				.b3(W2S103),
				.b4(W2S113),
				.b5(W2S123),
				.b6(W2S203),
				.b7(W2S213),
				.b8(W2S223),
				.c(c2312S)
);

ninexnine_unit ninexnine_unit_7080(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2S004),
				.b1(W2S014),
				.b2(W2S024),
				.b3(W2S104),
				.b4(W2S114),
				.b5(W2S124),
				.b6(W2S204),
				.b7(W2S214),
				.b8(W2S224),
				.c(c2412S)
);

ninexnine_unit ninexnine_unit_7081(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2S005),
				.b1(W2S015),
				.b2(W2S025),
				.b3(W2S105),
				.b4(W2S115),
				.b5(W2S125),
				.b6(W2S205),
				.b7(W2S215),
				.b8(W2S225),
				.c(c2512S)
);

ninexnine_unit ninexnine_unit_7082(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2S006),
				.b1(W2S016),
				.b2(W2S026),
				.b3(W2S106),
				.b4(W2S116),
				.b5(W2S126),
				.b6(W2S206),
				.b7(W2S216),
				.b8(W2S226),
				.c(c2612S)
);

ninexnine_unit ninexnine_unit_7083(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2S007),
				.b1(W2S017),
				.b2(W2S027),
				.b3(W2S107),
				.b4(W2S117),
				.b5(W2S127),
				.b6(W2S207),
				.b7(W2S217),
				.b8(W2S227),
				.c(c2712S)
);

ninexnine_unit ninexnine_unit_7084(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2S008),
				.b1(W2S018),
				.b2(W2S028),
				.b3(W2S108),
				.b4(W2S118),
				.b5(W2S128),
				.b6(W2S208),
				.b7(W2S218),
				.b8(W2S228),
				.c(c2812S)
);

ninexnine_unit ninexnine_unit_7085(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2S009),
				.b1(W2S019),
				.b2(W2S029),
				.b3(W2S109),
				.b4(W2S119),
				.b5(W2S129),
				.b6(W2S209),
				.b7(W2S219),
				.b8(W2S229),
				.c(c2912S)
);

ninexnine_unit ninexnine_unit_7086(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2S00A),
				.b1(W2S01A),
				.b2(W2S02A),
				.b3(W2S10A),
				.b4(W2S11A),
				.b5(W2S12A),
				.b6(W2S20A),
				.b7(W2S21A),
				.b8(W2S22A),
				.c(c2A12S)
);

ninexnine_unit ninexnine_unit_7087(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2S00B),
				.b1(W2S01B),
				.b2(W2S02B),
				.b3(W2S10B),
				.b4(W2S11B),
				.b5(W2S12B),
				.b6(W2S20B),
				.b7(W2S21B),
				.b8(W2S22B),
				.c(c2B12S)
);

ninexnine_unit ninexnine_unit_7088(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2S00C),
				.b1(W2S01C),
				.b2(W2S02C),
				.b3(W2S10C),
				.b4(W2S11C),
				.b5(W2S12C),
				.b6(W2S20C),
				.b7(W2S21C),
				.b8(W2S22C),
				.c(c2C12S)
);

ninexnine_unit ninexnine_unit_7089(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2S00D),
				.b1(W2S01D),
				.b2(W2S02D),
				.b3(W2S10D),
				.b4(W2S11D),
				.b5(W2S12D),
				.b6(W2S20D),
				.b7(W2S21D),
				.b8(W2S22D),
				.c(c2D12S)
);

ninexnine_unit ninexnine_unit_7090(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2S00E),
				.b1(W2S01E),
				.b2(W2S02E),
				.b3(W2S10E),
				.b4(W2S11E),
				.b5(W2S12E),
				.b6(W2S20E),
				.b7(W2S21E),
				.b8(W2S22E),
				.c(c2E12S)
);

ninexnine_unit ninexnine_unit_7091(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2S00F),
				.b1(W2S01F),
				.b2(W2S02F),
				.b3(W2S10F),
				.b4(W2S11F),
				.b5(W2S12F),
				.b6(W2S20F),
				.b7(W2S21F),
				.b8(W2S22F),
				.c(c2F12S)
);

assign C212S=c2012S+c2112S+c2212S+c2312S+c2412S+c2512S+c2612S+c2712S+c2812S+c2912S+c2A12S+c2B12S+c2C12S+c2D12S+c2E12S+c2F12S;
assign A212S=(C212S>=0)?1:0;

assign P312S=A212S;

ninexnine_unit ninexnine_unit_7092(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2S000),
				.b1(W2S010),
				.b2(W2S020),
				.b3(W2S100),
				.b4(W2S110),
				.b5(W2S120),
				.b6(W2S200),
				.b7(W2S210),
				.b8(W2S220),
				.c(c2020S)
);

ninexnine_unit ninexnine_unit_7093(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2S001),
				.b1(W2S011),
				.b2(W2S021),
				.b3(W2S101),
				.b4(W2S111),
				.b5(W2S121),
				.b6(W2S201),
				.b7(W2S211),
				.b8(W2S221),
				.c(c2120S)
);

ninexnine_unit ninexnine_unit_7094(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2S002),
				.b1(W2S012),
				.b2(W2S022),
				.b3(W2S102),
				.b4(W2S112),
				.b5(W2S122),
				.b6(W2S202),
				.b7(W2S212),
				.b8(W2S222),
				.c(c2220S)
);

ninexnine_unit ninexnine_unit_7095(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2S003),
				.b1(W2S013),
				.b2(W2S023),
				.b3(W2S103),
				.b4(W2S113),
				.b5(W2S123),
				.b6(W2S203),
				.b7(W2S213),
				.b8(W2S223),
				.c(c2320S)
);

ninexnine_unit ninexnine_unit_7096(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2S004),
				.b1(W2S014),
				.b2(W2S024),
				.b3(W2S104),
				.b4(W2S114),
				.b5(W2S124),
				.b6(W2S204),
				.b7(W2S214),
				.b8(W2S224),
				.c(c2420S)
);

ninexnine_unit ninexnine_unit_7097(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2S005),
				.b1(W2S015),
				.b2(W2S025),
				.b3(W2S105),
				.b4(W2S115),
				.b5(W2S125),
				.b6(W2S205),
				.b7(W2S215),
				.b8(W2S225),
				.c(c2520S)
);

ninexnine_unit ninexnine_unit_7098(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2S006),
				.b1(W2S016),
				.b2(W2S026),
				.b3(W2S106),
				.b4(W2S116),
				.b5(W2S126),
				.b6(W2S206),
				.b7(W2S216),
				.b8(W2S226),
				.c(c2620S)
);

ninexnine_unit ninexnine_unit_7099(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2S007),
				.b1(W2S017),
				.b2(W2S027),
				.b3(W2S107),
				.b4(W2S117),
				.b5(W2S127),
				.b6(W2S207),
				.b7(W2S217),
				.b8(W2S227),
				.c(c2720S)
);

ninexnine_unit ninexnine_unit_7100(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2S008),
				.b1(W2S018),
				.b2(W2S028),
				.b3(W2S108),
				.b4(W2S118),
				.b5(W2S128),
				.b6(W2S208),
				.b7(W2S218),
				.b8(W2S228),
				.c(c2820S)
);

ninexnine_unit ninexnine_unit_7101(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2S009),
				.b1(W2S019),
				.b2(W2S029),
				.b3(W2S109),
				.b4(W2S119),
				.b5(W2S129),
				.b6(W2S209),
				.b7(W2S219),
				.b8(W2S229),
				.c(c2920S)
);

ninexnine_unit ninexnine_unit_7102(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2S00A),
				.b1(W2S01A),
				.b2(W2S02A),
				.b3(W2S10A),
				.b4(W2S11A),
				.b5(W2S12A),
				.b6(W2S20A),
				.b7(W2S21A),
				.b8(W2S22A),
				.c(c2A20S)
);

ninexnine_unit ninexnine_unit_7103(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2S00B),
				.b1(W2S01B),
				.b2(W2S02B),
				.b3(W2S10B),
				.b4(W2S11B),
				.b5(W2S12B),
				.b6(W2S20B),
				.b7(W2S21B),
				.b8(W2S22B),
				.c(c2B20S)
);

ninexnine_unit ninexnine_unit_7104(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2S00C),
				.b1(W2S01C),
				.b2(W2S02C),
				.b3(W2S10C),
				.b4(W2S11C),
				.b5(W2S12C),
				.b6(W2S20C),
				.b7(W2S21C),
				.b8(W2S22C),
				.c(c2C20S)
);

ninexnine_unit ninexnine_unit_7105(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2S00D),
				.b1(W2S01D),
				.b2(W2S02D),
				.b3(W2S10D),
				.b4(W2S11D),
				.b5(W2S12D),
				.b6(W2S20D),
				.b7(W2S21D),
				.b8(W2S22D),
				.c(c2D20S)
);

ninexnine_unit ninexnine_unit_7106(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2S00E),
				.b1(W2S01E),
				.b2(W2S02E),
				.b3(W2S10E),
				.b4(W2S11E),
				.b5(W2S12E),
				.b6(W2S20E),
				.b7(W2S21E),
				.b8(W2S22E),
				.c(c2E20S)
);

ninexnine_unit ninexnine_unit_7107(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2S00F),
				.b1(W2S01F),
				.b2(W2S02F),
				.b3(W2S10F),
				.b4(W2S11F),
				.b5(W2S12F),
				.b6(W2S20F),
				.b7(W2S21F),
				.b8(W2S22F),
				.c(c2F20S)
);

assign C220S=c2020S+c2120S+c2220S+c2320S+c2420S+c2520S+c2620S+c2720S+c2820S+c2920S+c2A20S+c2B20S+c2C20S+c2D20S+c2E20S+c2F20S;
assign A220S=(C220S>=0)?1:0;

assign P320S=A220S;

ninexnine_unit ninexnine_unit_7108(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2S000),
				.b1(W2S010),
				.b2(W2S020),
				.b3(W2S100),
				.b4(W2S110),
				.b5(W2S120),
				.b6(W2S200),
				.b7(W2S210),
				.b8(W2S220),
				.c(c2021S)
);

ninexnine_unit ninexnine_unit_7109(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2S001),
				.b1(W2S011),
				.b2(W2S021),
				.b3(W2S101),
				.b4(W2S111),
				.b5(W2S121),
				.b6(W2S201),
				.b7(W2S211),
				.b8(W2S221),
				.c(c2121S)
);

ninexnine_unit ninexnine_unit_7110(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2S002),
				.b1(W2S012),
				.b2(W2S022),
				.b3(W2S102),
				.b4(W2S112),
				.b5(W2S122),
				.b6(W2S202),
				.b7(W2S212),
				.b8(W2S222),
				.c(c2221S)
);

ninexnine_unit ninexnine_unit_7111(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2S003),
				.b1(W2S013),
				.b2(W2S023),
				.b3(W2S103),
				.b4(W2S113),
				.b5(W2S123),
				.b6(W2S203),
				.b7(W2S213),
				.b8(W2S223),
				.c(c2321S)
);

ninexnine_unit ninexnine_unit_7112(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2S004),
				.b1(W2S014),
				.b2(W2S024),
				.b3(W2S104),
				.b4(W2S114),
				.b5(W2S124),
				.b6(W2S204),
				.b7(W2S214),
				.b8(W2S224),
				.c(c2421S)
);

ninexnine_unit ninexnine_unit_7113(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2S005),
				.b1(W2S015),
				.b2(W2S025),
				.b3(W2S105),
				.b4(W2S115),
				.b5(W2S125),
				.b6(W2S205),
				.b7(W2S215),
				.b8(W2S225),
				.c(c2521S)
);

ninexnine_unit ninexnine_unit_7114(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2S006),
				.b1(W2S016),
				.b2(W2S026),
				.b3(W2S106),
				.b4(W2S116),
				.b5(W2S126),
				.b6(W2S206),
				.b7(W2S216),
				.b8(W2S226),
				.c(c2621S)
);

ninexnine_unit ninexnine_unit_7115(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2S007),
				.b1(W2S017),
				.b2(W2S027),
				.b3(W2S107),
				.b4(W2S117),
				.b5(W2S127),
				.b6(W2S207),
				.b7(W2S217),
				.b8(W2S227),
				.c(c2721S)
);

ninexnine_unit ninexnine_unit_7116(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2S008),
				.b1(W2S018),
				.b2(W2S028),
				.b3(W2S108),
				.b4(W2S118),
				.b5(W2S128),
				.b6(W2S208),
				.b7(W2S218),
				.b8(W2S228),
				.c(c2821S)
);

ninexnine_unit ninexnine_unit_7117(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2S009),
				.b1(W2S019),
				.b2(W2S029),
				.b3(W2S109),
				.b4(W2S119),
				.b5(W2S129),
				.b6(W2S209),
				.b7(W2S219),
				.b8(W2S229),
				.c(c2921S)
);

ninexnine_unit ninexnine_unit_7118(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2S00A),
				.b1(W2S01A),
				.b2(W2S02A),
				.b3(W2S10A),
				.b4(W2S11A),
				.b5(W2S12A),
				.b6(W2S20A),
				.b7(W2S21A),
				.b8(W2S22A),
				.c(c2A21S)
);

ninexnine_unit ninexnine_unit_7119(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2S00B),
				.b1(W2S01B),
				.b2(W2S02B),
				.b3(W2S10B),
				.b4(W2S11B),
				.b5(W2S12B),
				.b6(W2S20B),
				.b7(W2S21B),
				.b8(W2S22B),
				.c(c2B21S)
);

ninexnine_unit ninexnine_unit_7120(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2S00C),
				.b1(W2S01C),
				.b2(W2S02C),
				.b3(W2S10C),
				.b4(W2S11C),
				.b5(W2S12C),
				.b6(W2S20C),
				.b7(W2S21C),
				.b8(W2S22C),
				.c(c2C21S)
);

ninexnine_unit ninexnine_unit_7121(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2S00D),
				.b1(W2S01D),
				.b2(W2S02D),
				.b3(W2S10D),
				.b4(W2S11D),
				.b5(W2S12D),
				.b6(W2S20D),
				.b7(W2S21D),
				.b8(W2S22D),
				.c(c2D21S)
);

ninexnine_unit ninexnine_unit_7122(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2S00E),
				.b1(W2S01E),
				.b2(W2S02E),
				.b3(W2S10E),
				.b4(W2S11E),
				.b5(W2S12E),
				.b6(W2S20E),
				.b7(W2S21E),
				.b8(W2S22E),
				.c(c2E21S)
);

ninexnine_unit ninexnine_unit_7123(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2S00F),
				.b1(W2S01F),
				.b2(W2S02F),
				.b3(W2S10F),
				.b4(W2S11F),
				.b5(W2S12F),
				.b6(W2S20F),
				.b7(W2S21F),
				.b8(W2S22F),
				.c(c2F21S)
);

assign C221S=c2021S+c2121S+c2221S+c2321S+c2421S+c2521S+c2621S+c2721S+c2821S+c2921S+c2A21S+c2B21S+c2C21S+c2D21S+c2E21S+c2F21S;
assign A221S=(C221S>=0)?1:0;

assign P321S=A221S;

ninexnine_unit ninexnine_unit_7124(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2S000),
				.b1(W2S010),
				.b2(W2S020),
				.b3(W2S100),
				.b4(W2S110),
				.b5(W2S120),
				.b6(W2S200),
				.b7(W2S210),
				.b8(W2S220),
				.c(c2022S)
);

ninexnine_unit ninexnine_unit_7125(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2S001),
				.b1(W2S011),
				.b2(W2S021),
				.b3(W2S101),
				.b4(W2S111),
				.b5(W2S121),
				.b6(W2S201),
				.b7(W2S211),
				.b8(W2S221),
				.c(c2122S)
);

ninexnine_unit ninexnine_unit_7126(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2S002),
				.b1(W2S012),
				.b2(W2S022),
				.b3(W2S102),
				.b4(W2S112),
				.b5(W2S122),
				.b6(W2S202),
				.b7(W2S212),
				.b8(W2S222),
				.c(c2222S)
);

ninexnine_unit ninexnine_unit_7127(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2S003),
				.b1(W2S013),
				.b2(W2S023),
				.b3(W2S103),
				.b4(W2S113),
				.b5(W2S123),
				.b6(W2S203),
				.b7(W2S213),
				.b8(W2S223),
				.c(c2322S)
);

ninexnine_unit ninexnine_unit_7128(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2S004),
				.b1(W2S014),
				.b2(W2S024),
				.b3(W2S104),
				.b4(W2S114),
				.b5(W2S124),
				.b6(W2S204),
				.b7(W2S214),
				.b8(W2S224),
				.c(c2422S)
);

ninexnine_unit ninexnine_unit_7129(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2S005),
				.b1(W2S015),
				.b2(W2S025),
				.b3(W2S105),
				.b4(W2S115),
				.b5(W2S125),
				.b6(W2S205),
				.b7(W2S215),
				.b8(W2S225),
				.c(c2522S)
);

ninexnine_unit ninexnine_unit_7130(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2S006),
				.b1(W2S016),
				.b2(W2S026),
				.b3(W2S106),
				.b4(W2S116),
				.b5(W2S126),
				.b6(W2S206),
				.b7(W2S216),
				.b8(W2S226),
				.c(c2622S)
);

ninexnine_unit ninexnine_unit_7131(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2S007),
				.b1(W2S017),
				.b2(W2S027),
				.b3(W2S107),
				.b4(W2S117),
				.b5(W2S127),
				.b6(W2S207),
				.b7(W2S217),
				.b8(W2S227),
				.c(c2722S)
);

ninexnine_unit ninexnine_unit_7132(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2S008),
				.b1(W2S018),
				.b2(W2S028),
				.b3(W2S108),
				.b4(W2S118),
				.b5(W2S128),
				.b6(W2S208),
				.b7(W2S218),
				.b8(W2S228),
				.c(c2822S)
);

ninexnine_unit ninexnine_unit_7133(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2S009),
				.b1(W2S019),
				.b2(W2S029),
				.b3(W2S109),
				.b4(W2S119),
				.b5(W2S129),
				.b6(W2S209),
				.b7(W2S219),
				.b8(W2S229),
				.c(c2922S)
);

ninexnine_unit ninexnine_unit_7134(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2S00A),
				.b1(W2S01A),
				.b2(W2S02A),
				.b3(W2S10A),
				.b4(W2S11A),
				.b5(W2S12A),
				.b6(W2S20A),
				.b7(W2S21A),
				.b8(W2S22A),
				.c(c2A22S)
);

ninexnine_unit ninexnine_unit_7135(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2S00B),
				.b1(W2S01B),
				.b2(W2S02B),
				.b3(W2S10B),
				.b4(W2S11B),
				.b5(W2S12B),
				.b6(W2S20B),
				.b7(W2S21B),
				.b8(W2S22B),
				.c(c2B22S)
);

ninexnine_unit ninexnine_unit_7136(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2S00C),
				.b1(W2S01C),
				.b2(W2S02C),
				.b3(W2S10C),
				.b4(W2S11C),
				.b5(W2S12C),
				.b6(W2S20C),
				.b7(W2S21C),
				.b8(W2S22C),
				.c(c2C22S)
);

ninexnine_unit ninexnine_unit_7137(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2S00D),
				.b1(W2S01D),
				.b2(W2S02D),
				.b3(W2S10D),
				.b4(W2S11D),
				.b5(W2S12D),
				.b6(W2S20D),
				.b7(W2S21D),
				.b8(W2S22D),
				.c(c2D22S)
);

ninexnine_unit ninexnine_unit_7138(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2S00E),
				.b1(W2S01E),
				.b2(W2S02E),
				.b3(W2S10E),
				.b4(W2S11E),
				.b5(W2S12E),
				.b6(W2S20E),
				.b7(W2S21E),
				.b8(W2S22E),
				.c(c2E22S)
);

ninexnine_unit ninexnine_unit_7139(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2S00F),
				.b1(W2S01F),
				.b2(W2S02F),
				.b3(W2S10F),
				.b4(W2S11F),
				.b5(W2S12F),
				.b6(W2S20F),
				.b7(W2S21F),
				.b8(W2S22F),
				.c(c2F22S)
);

assign C222S=c2022S+c2122S+c2222S+c2322S+c2422S+c2522S+c2622S+c2722S+c2822S+c2922S+c2A22S+c2B22S+c2C22S+c2D22S+c2E22S+c2F22S;
assign A222S=(C222S>=0)?1:0;

assign P322S=A222S;

ninexnine_unit ninexnine_unit_7140(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2T000),
				.b1(W2T010),
				.b2(W2T020),
				.b3(W2T100),
				.b4(W2T110),
				.b5(W2T120),
				.b6(W2T200),
				.b7(W2T210),
				.b8(W2T220),
				.c(c2000T)
);

ninexnine_unit ninexnine_unit_7141(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2T001),
				.b1(W2T011),
				.b2(W2T021),
				.b3(W2T101),
				.b4(W2T111),
				.b5(W2T121),
				.b6(W2T201),
				.b7(W2T211),
				.b8(W2T221),
				.c(c2100T)
);

ninexnine_unit ninexnine_unit_7142(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2T002),
				.b1(W2T012),
				.b2(W2T022),
				.b3(W2T102),
				.b4(W2T112),
				.b5(W2T122),
				.b6(W2T202),
				.b7(W2T212),
				.b8(W2T222),
				.c(c2200T)
);

ninexnine_unit ninexnine_unit_7143(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2T003),
				.b1(W2T013),
				.b2(W2T023),
				.b3(W2T103),
				.b4(W2T113),
				.b5(W2T123),
				.b6(W2T203),
				.b7(W2T213),
				.b8(W2T223),
				.c(c2300T)
);

ninexnine_unit ninexnine_unit_7144(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2T004),
				.b1(W2T014),
				.b2(W2T024),
				.b3(W2T104),
				.b4(W2T114),
				.b5(W2T124),
				.b6(W2T204),
				.b7(W2T214),
				.b8(W2T224),
				.c(c2400T)
);

ninexnine_unit ninexnine_unit_7145(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2T005),
				.b1(W2T015),
				.b2(W2T025),
				.b3(W2T105),
				.b4(W2T115),
				.b5(W2T125),
				.b6(W2T205),
				.b7(W2T215),
				.b8(W2T225),
				.c(c2500T)
);

ninexnine_unit ninexnine_unit_7146(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2T006),
				.b1(W2T016),
				.b2(W2T026),
				.b3(W2T106),
				.b4(W2T116),
				.b5(W2T126),
				.b6(W2T206),
				.b7(W2T216),
				.b8(W2T226),
				.c(c2600T)
);

ninexnine_unit ninexnine_unit_7147(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2T007),
				.b1(W2T017),
				.b2(W2T027),
				.b3(W2T107),
				.b4(W2T117),
				.b5(W2T127),
				.b6(W2T207),
				.b7(W2T217),
				.b8(W2T227),
				.c(c2700T)
);

ninexnine_unit ninexnine_unit_7148(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2T008),
				.b1(W2T018),
				.b2(W2T028),
				.b3(W2T108),
				.b4(W2T118),
				.b5(W2T128),
				.b6(W2T208),
				.b7(W2T218),
				.b8(W2T228),
				.c(c2800T)
);

ninexnine_unit ninexnine_unit_7149(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2T009),
				.b1(W2T019),
				.b2(W2T029),
				.b3(W2T109),
				.b4(W2T119),
				.b5(W2T129),
				.b6(W2T209),
				.b7(W2T219),
				.b8(W2T229),
				.c(c2900T)
);

ninexnine_unit ninexnine_unit_7150(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2T00A),
				.b1(W2T01A),
				.b2(W2T02A),
				.b3(W2T10A),
				.b4(W2T11A),
				.b5(W2T12A),
				.b6(W2T20A),
				.b7(W2T21A),
				.b8(W2T22A),
				.c(c2A00T)
);

ninexnine_unit ninexnine_unit_7151(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2T00B),
				.b1(W2T01B),
				.b2(W2T02B),
				.b3(W2T10B),
				.b4(W2T11B),
				.b5(W2T12B),
				.b6(W2T20B),
				.b7(W2T21B),
				.b8(W2T22B),
				.c(c2B00T)
);

ninexnine_unit ninexnine_unit_7152(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2T00C),
				.b1(W2T01C),
				.b2(W2T02C),
				.b3(W2T10C),
				.b4(W2T11C),
				.b5(W2T12C),
				.b6(W2T20C),
				.b7(W2T21C),
				.b8(W2T22C),
				.c(c2C00T)
);

ninexnine_unit ninexnine_unit_7153(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2T00D),
				.b1(W2T01D),
				.b2(W2T02D),
				.b3(W2T10D),
				.b4(W2T11D),
				.b5(W2T12D),
				.b6(W2T20D),
				.b7(W2T21D),
				.b8(W2T22D),
				.c(c2D00T)
);

ninexnine_unit ninexnine_unit_7154(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2T00E),
				.b1(W2T01E),
				.b2(W2T02E),
				.b3(W2T10E),
				.b4(W2T11E),
				.b5(W2T12E),
				.b6(W2T20E),
				.b7(W2T21E),
				.b8(W2T22E),
				.c(c2E00T)
);

ninexnine_unit ninexnine_unit_7155(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2T00F),
				.b1(W2T01F),
				.b2(W2T02F),
				.b3(W2T10F),
				.b4(W2T11F),
				.b5(W2T12F),
				.b6(W2T20F),
				.b7(W2T21F),
				.b8(W2T22F),
				.c(c2F00T)
);

assign C200T=c2000T+c2100T+c2200T+c2300T+c2400T+c2500T+c2600T+c2700T+c2800T+c2900T+c2A00T+c2B00T+c2C00T+c2D00T+c2E00T+c2F00T;
assign A200T=(C200T>=0)?1:0;

assign P300T=A200T;

ninexnine_unit ninexnine_unit_7156(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2T000),
				.b1(W2T010),
				.b2(W2T020),
				.b3(W2T100),
				.b4(W2T110),
				.b5(W2T120),
				.b6(W2T200),
				.b7(W2T210),
				.b8(W2T220),
				.c(c2001T)
);

ninexnine_unit ninexnine_unit_7157(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2T001),
				.b1(W2T011),
				.b2(W2T021),
				.b3(W2T101),
				.b4(W2T111),
				.b5(W2T121),
				.b6(W2T201),
				.b7(W2T211),
				.b8(W2T221),
				.c(c2101T)
);

ninexnine_unit ninexnine_unit_7158(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2T002),
				.b1(W2T012),
				.b2(W2T022),
				.b3(W2T102),
				.b4(W2T112),
				.b5(W2T122),
				.b6(W2T202),
				.b7(W2T212),
				.b8(W2T222),
				.c(c2201T)
);

ninexnine_unit ninexnine_unit_7159(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2T003),
				.b1(W2T013),
				.b2(W2T023),
				.b3(W2T103),
				.b4(W2T113),
				.b5(W2T123),
				.b6(W2T203),
				.b7(W2T213),
				.b8(W2T223),
				.c(c2301T)
);

ninexnine_unit ninexnine_unit_7160(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2T004),
				.b1(W2T014),
				.b2(W2T024),
				.b3(W2T104),
				.b4(W2T114),
				.b5(W2T124),
				.b6(W2T204),
				.b7(W2T214),
				.b8(W2T224),
				.c(c2401T)
);

ninexnine_unit ninexnine_unit_7161(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2T005),
				.b1(W2T015),
				.b2(W2T025),
				.b3(W2T105),
				.b4(W2T115),
				.b5(W2T125),
				.b6(W2T205),
				.b7(W2T215),
				.b8(W2T225),
				.c(c2501T)
);

ninexnine_unit ninexnine_unit_7162(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2T006),
				.b1(W2T016),
				.b2(W2T026),
				.b3(W2T106),
				.b4(W2T116),
				.b5(W2T126),
				.b6(W2T206),
				.b7(W2T216),
				.b8(W2T226),
				.c(c2601T)
);

ninexnine_unit ninexnine_unit_7163(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2T007),
				.b1(W2T017),
				.b2(W2T027),
				.b3(W2T107),
				.b4(W2T117),
				.b5(W2T127),
				.b6(W2T207),
				.b7(W2T217),
				.b8(W2T227),
				.c(c2701T)
);

ninexnine_unit ninexnine_unit_7164(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2T008),
				.b1(W2T018),
				.b2(W2T028),
				.b3(W2T108),
				.b4(W2T118),
				.b5(W2T128),
				.b6(W2T208),
				.b7(W2T218),
				.b8(W2T228),
				.c(c2801T)
);

ninexnine_unit ninexnine_unit_7165(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2T009),
				.b1(W2T019),
				.b2(W2T029),
				.b3(W2T109),
				.b4(W2T119),
				.b5(W2T129),
				.b6(W2T209),
				.b7(W2T219),
				.b8(W2T229),
				.c(c2901T)
);

ninexnine_unit ninexnine_unit_7166(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2T00A),
				.b1(W2T01A),
				.b2(W2T02A),
				.b3(W2T10A),
				.b4(W2T11A),
				.b5(W2T12A),
				.b6(W2T20A),
				.b7(W2T21A),
				.b8(W2T22A),
				.c(c2A01T)
);

ninexnine_unit ninexnine_unit_7167(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2T00B),
				.b1(W2T01B),
				.b2(W2T02B),
				.b3(W2T10B),
				.b4(W2T11B),
				.b5(W2T12B),
				.b6(W2T20B),
				.b7(W2T21B),
				.b8(W2T22B),
				.c(c2B01T)
);

ninexnine_unit ninexnine_unit_7168(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2T00C),
				.b1(W2T01C),
				.b2(W2T02C),
				.b3(W2T10C),
				.b4(W2T11C),
				.b5(W2T12C),
				.b6(W2T20C),
				.b7(W2T21C),
				.b8(W2T22C),
				.c(c2C01T)
);

ninexnine_unit ninexnine_unit_7169(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2T00D),
				.b1(W2T01D),
				.b2(W2T02D),
				.b3(W2T10D),
				.b4(W2T11D),
				.b5(W2T12D),
				.b6(W2T20D),
				.b7(W2T21D),
				.b8(W2T22D),
				.c(c2D01T)
);

ninexnine_unit ninexnine_unit_7170(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2T00E),
				.b1(W2T01E),
				.b2(W2T02E),
				.b3(W2T10E),
				.b4(W2T11E),
				.b5(W2T12E),
				.b6(W2T20E),
				.b7(W2T21E),
				.b8(W2T22E),
				.c(c2E01T)
);

ninexnine_unit ninexnine_unit_7171(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2T00F),
				.b1(W2T01F),
				.b2(W2T02F),
				.b3(W2T10F),
				.b4(W2T11F),
				.b5(W2T12F),
				.b6(W2T20F),
				.b7(W2T21F),
				.b8(W2T22F),
				.c(c2F01T)
);

assign C201T=c2001T+c2101T+c2201T+c2301T+c2401T+c2501T+c2601T+c2701T+c2801T+c2901T+c2A01T+c2B01T+c2C01T+c2D01T+c2E01T+c2F01T;
assign A201T=(C201T>=0)?1:0;

assign P301T=A201T;

ninexnine_unit ninexnine_unit_7172(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2T000),
				.b1(W2T010),
				.b2(W2T020),
				.b3(W2T100),
				.b4(W2T110),
				.b5(W2T120),
				.b6(W2T200),
				.b7(W2T210),
				.b8(W2T220),
				.c(c2002T)
);

ninexnine_unit ninexnine_unit_7173(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2T001),
				.b1(W2T011),
				.b2(W2T021),
				.b3(W2T101),
				.b4(W2T111),
				.b5(W2T121),
				.b6(W2T201),
				.b7(W2T211),
				.b8(W2T221),
				.c(c2102T)
);

ninexnine_unit ninexnine_unit_7174(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2T002),
				.b1(W2T012),
				.b2(W2T022),
				.b3(W2T102),
				.b4(W2T112),
				.b5(W2T122),
				.b6(W2T202),
				.b7(W2T212),
				.b8(W2T222),
				.c(c2202T)
);

ninexnine_unit ninexnine_unit_7175(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2T003),
				.b1(W2T013),
				.b2(W2T023),
				.b3(W2T103),
				.b4(W2T113),
				.b5(W2T123),
				.b6(W2T203),
				.b7(W2T213),
				.b8(W2T223),
				.c(c2302T)
);

ninexnine_unit ninexnine_unit_7176(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2T004),
				.b1(W2T014),
				.b2(W2T024),
				.b3(W2T104),
				.b4(W2T114),
				.b5(W2T124),
				.b6(W2T204),
				.b7(W2T214),
				.b8(W2T224),
				.c(c2402T)
);

ninexnine_unit ninexnine_unit_7177(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2T005),
				.b1(W2T015),
				.b2(W2T025),
				.b3(W2T105),
				.b4(W2T115),
				.b5(W2T125),
				.b6(W2T205),
				.b7(W2T215),
				.b8(W2T225),
				.c(c2502T)
);

ninexnine_unit ninexnine_unit_7178(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2T006),
				.b1(W2T016),
				.b2(W2T026),
				.b3(W2T106),
				.b4(W2T116),
				.b5(W2T126),
				.b6(W2T206),
				.b7(W2T216),
				.b8(W2T226),
				.c(c2602T)
);

ninexnine_unit ninexnine_unit_7179(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2T007),
				.b1(W2T017),
				.b2(W2T027),
				.b3(W2T107),
				.b4(W2T117),
				.b5(W2T127),
				.b6(W2T207),
				.b7(W2T217),
				.b8(W2T227),
				.c(c2702T)
);

ninexnine_unit ninexnine_unit_7180(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2T008),
				.b1(W2T018),
				.b2(W2T028),
				.b3(W2T108),
				.b4(W2T118),
				.b5(W2T128),
				.b6(W2T208),
				.b7(W2T218),
				.b8(W2T228),
				.c(c2802T)
);

ninexnine_unit ninexnine_unit_7181(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2T009),
				.b1(W2T019),
				.b2(W2T029),
				.b3(W2T109),
				.b4(W2T119),
				.b5(W2T129),
				.b6(W2T209),
				.b7(W2T219),
				.b8(W2T229),
				.c(c2902T)
);

ninexnine_unit ninexnine_unit_7182(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2T00A),
				.b1(W2T01A),
				.b2(W2T02A),
				.b3(W2T10A),
				.b4(W2T11A),
				.b5(W2T12A),
				.b6(W2T20A),
				.b7(W2T21A),
				.b8(W2T22A),
				.c(c2A02T)
);

ninexnine_unit ninexnine_unit_7183(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2T00B),
				.b1(W2T01B),
				.b2(W2T02B),
				.b3(W2T10B),
				.b4(W2T11B),
				.b5(W2T12B),
				.b6(W2T20B),
				.b7(W2T21B),
				.b8(W2T22B),
				.c(c2B02T)
);

ninexnine_unit ninexnine_unit_7184(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2T00C),
				.b1(W2T01C),
				.b2(W2T02C),
				.b3(W2T10C),
				.b4(W2T11C),
				.b5(W2T12C),
				.b6(W2T20C),
				.b7(W2T21C),
				.b8(W2T22C),
				.c(c2C02T)
);

ninexnine_unit ninexnine_unit_7185(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2T00D),
				.b1(W2T01D),
				.b2(W2T02D),
				.b3(W2T10D),
				.b4(W2T11D),
				.b5(W2T12D),
				.b6(W2T20D),
				.b7(W2T21D),
				.b8(W2T22D),
				.c(c2D02T)
);

ninexnine_unit ninexnine_unit_7186(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2T00E),
				.b1(W2T01E),
				.b2(W2T02E),
				.b3(W2T10E),
				.b4(W2T11E),
				.b5(W2T12E),
				.b6(W2T20E),
				.b7(W2T21E),
				.b8(W2T22E),
				.c(c2E02T)
);

ninexnine_unit ninexnine_unit_7187(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2T00F),
				.b1(W2T01F),
				.b2(W2T02F),
				.b3(W2T10F),
				.b4(W2T11F),
				.b5(W2T12F),
				.b6(W2T20F),
				.b7(W2T21F),
				.b8(W2T22F),
				.c(c2F02T)
);

assign C202T=c2002T+c2102T+c2202T+c2302T+c2402T+c2502T+c2602T+c2702T+c2802T+c2902T+c2A02T+c2B02T+c2C02T+c2D02T+c2E02T+c2F02T;
assign A202T=(C202T>=0)?1:0;

assign P302T=A202T;

ninexnine_unit ninexnine_unit_7188(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2T000),
				.b1(W2T010),
				.b2(W2T020),
				.b3(W2T100),
				.b4(W2T110),
				.b5(W2T120),
				.b6(W2T200),
				.b7(W2T210),
				.b8(W2T220),
				.c(c2010T)
);

ninexnine_unit ninexnine_unit_7189(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2T001),
				.b1(W2T011),
				.b2(W2T021),
				.b3(W2T101),
				.b4(W2T111),
				.b5(W2T121),
				.b6(W2T201),
				.b7(W2T211),
				.b8(W2T221),
				.c(c2110T)
);

ninexnine_unit ninexnine_unit_7190(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2T002),
				.b1(W2T012),
				.b2(W2T022),
				.b3(W2T102),
				.b4(W2T112),
				.b5(W2T122),
				.b6(W2T202),
				.b7(W2T212),
				.b8(W2T222),
				.c(c2210T)
);

ninexnine_unit ninexnine_unit_7191(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2T003),
				.b1(W2T013),
				.b2(W2T023),
				.b3(W2T103),
				.b4(W2T113),
				.b5(W2T123),
				.b6(W2T203),
				.b7(W2T213),
				.b8(W2T223),
				.c(c2310T)
);

ninexnine_unit ninexnine_unit_7192(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2T004),
				.b1(W2T014),
				.b2(W2T024),
				.b3(W2T104),
				.b4(W2T114),
				.b5(W2T124),
				.b6(W2T204),
				.b7(W2T214),
				.b8(W2T224),
				.c(c2410T)
);

ninexnine_unit ninexnine_unit_7193(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2T005),
				.b1(W2T015),
				.b2(W2T025),
				.b3(W2T105),
				.b4(W2T115),
				.b5(W2T125),
				.b6(W2T205),
				.b7(W2T215),
				.b8(W2T225),
				.c(c2510T)
);

ninexnine_unit ninexnine_unit_7194(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2T006),
				.b1(W2T016),
				.b2(W2T026),
				.b3(W2T106),
				.b4(W2T116),
				.b5(W2T126),
				.b6(W2T206),
				.b7(W2T216),
				.b8(W2T226),
				.c(c2610T)
);

ninexnine_unit ninexnine_unit_7195(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2T007),
				.b1(W2T017),
				.b2(W2T027),
				.b3(W2T107),
				.b4(W2T117),
				.b5(W2T127),
				.b6(W2T207),
				.b7(W2T217),
				.b8(W2T227),
				.c(c2710T)
);

ninexnine_unit ninexnine_unit_7196(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2T008),
				.b1(W2T018),
				.b2(W2T028),
				.b3(W2T108),
				.b4(W2T118),
				.b5(W2T128),
				.b6(W2T208),
				.b7(W2T218),
				.b8(W2T228),
				.c(c2810T)
);

ninexnine_unit ninexnine_unit_7197(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2T009),
				.b1(W2T019),
				.b2(W2T029),
				.b3(W2T109),
				.b4(W2T119),
				.b5(W2T129),
				.b6(W2T209),
				.b7(W2T219),
				.b8(W2T229),
				.c(c2910T)
);

ninexnine_unit ninexnine_unit_7198(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2T00A),
				.b1(W2T01A),
				.b2(W2T02A),
				.b3(W2T10A),
				.b4(W2T11A),
				.b5(W2T12A),
				.b6(W2T20A),
				.b7(W2T21A),
				.b8(W2T22A),
				.c(c2A10T)
);

ninexnine_unit ninexnine_unit_7199(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2T00B),
				.b1(W2T01B),
				.b2(W2T02B),
				.b3(W2T10B),
				.b4(W2T11B),
				.b5(W2T12B),
				.b6(W2T20B),
				.b7(W2T21B),
				.b8(W2T22B),
				.c(c2B10T)
);

ninexnine_unit ninexnine_unit_7200(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2T00C),
				.b1(W2T01C),
				.b2(W2T02C),
				.b3(W2T10C),
				.b4(W2T11C),
				.b5(W2T12C),
				.b6(W2T20C),
				.b7(W2T21C),
				.b8(W2T22C),
				.c(c2C10T)
);

ninexnine_unit ninexnine_unit_7201(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2T00D),
				.b1(W2T01D),
				.b2(W2T02D),
				.b3(W2T10D),
				.b4(W2T11D),
				.b5(W2T12D),
				.b6(W2T20D),
				.b7(W2T21D),
				.b8(W2T22D),
				.c(c2D10T)
);

ninexnine_unit ninexnine_unit_7202(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2T00E),
				.b1(W2T01E),
				.b2(W2T02E),
				.b3(W2T10E),
				.b4(W2T11E),
				.b5(W2T12E),
				.b6(W2T20E),
				.b7(W2T21E),
				.b8(W2T22E),
				.c(c2E10T)
);

ninexnine_unit ninexnine_unit_7203(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2T00F),
				.b1(W2T01F),
				.b2(W2T02F),
				.b3(W2T10F),
				.b4(W2T11F),
				.b5(W2T12F),
				.b6(W2T20F),
				.b7(W2T21F),
				.b8(W2T22F),
				.c(c2F10T)
);

assign C210T=c2010T+c2110T+c2210T+c2310T+c2410T+c2510T+c2610T+c2710T+c2810T+c2910T+c2A10T+c2B10T+c2C10T+c2D10T+c2E10T+c2F10T;
assign A210T=(C210T>=0)?1:0;

assign P310T=A210T;

ninexnine_unit ninexnine_unit_7204(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2T000),
				.b1(W2T010),
				.b2(W2T020),
				.b3(W2T100),
				.b4(W2T110),
				.b5(W2T120),
				.b6(W2T200),
				.b7(W2T210),
				.b8(W2T220),
				.c(c2011T)
);

ninexnine_unit ninexnine_unit_7205(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2T001),
				.b1(W2T011),
				.b2(W2T021),
				.b3(W2T101),
				.b4(W2T111),
				.b5(W2T121),
				.b6(W2T201),
				.b7(W2T211),
				.b8(W2T221),
				.c(c2111T)
);

ninexnine_unit ninexnine_unit_7206(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2T002),
				.b1(W2T012),
				.b2(W2T022),
				.b3(W2T102),
				.b4(W2T112),
				.b5(W2T122),
				.b6(W2T202),
				.b7(W2T212),
				.b8(W2T222),
				.c(c2211T)
);

ninexnine_unit ninexnine_unit_7207(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2T003),
				.b1(W2T013),
				.b2(W2T023),
				.b3(W2T103),
				.b4(W2T113),
				.b5(W2T123),
				.b6(W2T203),
				.b7(W2T213),
				.b8(W2T223),
				.c(c2311T)
);

ninexnine_unit ninexnine_unit_7208(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2T004),
				.b1(W2T014),
				.b2(W2T024),
				.b3(W2T104),
				.b4(W2T114),
				.b5(W2T124),
				.b6(W2T204),
				.b7(W2T214),
				.b8(W2T224),
				.c(c2411T)
);

ninexnine_unit ninexnine_unit_7209(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2T005),
				.b1(W2T015),
				.b2(W2T025),
				.b3(W2T105),
				.b4(W2T115),
				.b5(W2T125),
				.b6(W2T205),
				.b7(W2T215),
				.b8(W2T225),
				.c(c2511T)
);

ninexnine_unit ninexnine_unit_7210(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2T006),
				.b1(W2T016),
				.b2(W2T026),
				.b3(W2T106),
				.b4(W2T116),
				.b5(W2T126),
				.b6(W2T206),
				.b7(W2T216),
				.b8(W2T226),
				.c(c2611T)
);

ninexnine_unit ninexnine_unit_7211(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2T007),
				.b1(W2T017),
				.b2(W2T027),
				.b3(W2T107),
				.b4(W2T117),
				.b5(W2T127),
				.b6(W2T207),
				.b7(W2T217),
				.b8(W2T227),
				.c(c2711T)
);

ninexnine_unit ninexnine_unit_7212(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2T008),
				.b1(W2T018),
				.b2(W2T028),
				.b3(W2T108),
				.b4(W2T118),
				.b5(W2T128),
				.b6(W2T208),
				.b7(W2T218),
				.b8(W2T228),
				.c(c2811T)
);

ninexnine_unit ninexnine_unit_7213(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2T009),
				.b1(W2T019),
				.b2(W2T029),
				.b3(W2T109),
				.b4(W2T119),
				.b5(W2T129),
				.b6(W2T209),
				.b7(W2T219),
				.b8(W2T229),
				.c(c2911T)
);

ninexnine_unit ninexnine_unit_7214(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2T00A),
				.b1(W2T01A),
				.b2(W2T02A),
				.b3(W2T10A),
				.b4(W2T11A),
				.b5(W2T12A),
				.b6(W2T20A),
				.b7(W2T21A),
				.b8(W2T22A),
				.c(c2A11T)
);

ninexnine_unit ninexnine_unit_7215(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2T00B),
				.b1(W2T01B),
				.b2(W2T02B),
				.b3(W2T10B),
				.b4(W2T11B),
				.b5(W2T12B),
				.b6(W2T20B),
				.b7(W2T21B),
				.b8(W2T22B),
				.c(c2B11T)
);

ninexnine_unit ninexnine_unit_7216(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2T00C),
				.b1(W2T01C),
				.b2(W2T02C),
				.b3(W2T10C),
				.b4(W2T11C),
				.b5(W2T12C),
				.b6(W2T20C),
				.b7(W2T21C),
				.b8(W2T22C),
				.c(c2C11T)
);

ninexnine_unit ninexnine_unit_7217(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2T00D),
				.b1(W2T01D),
				.b2(W2T02D),
				.b3(W2T10D),
				.b4(W2T11D),
				.b5(W2T12D),
				.b6(W2T20D),
				.b7(W2T21D),
				.b8(W2T22D),
				.c(c2D11T)
);

ninexnine_unit ninexnine_unit_7218(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2T00E),
				.b1(W2T01E),
				.b2(W2T02E),
				.b3(W2T10E),
				.b4(W2T11E),
				.b5(W2T12E),
				.b6(W2T20E),
				.b7(W2T21E),
				.b8(W2T22E),
				.c(c2E11T)
);

ninexnine_unit ninexnine_unit_7219(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2T00F),
				.b1(W2T01F),
				.b2(W2T02F),
				.b3(W2T10F),
				.b4(W2T11F),
				.b5(W2T12F),
				.b6(W2T20F),
				.b7(W2T21F),
				.b8(W2T22F),
				.c(c2F11T)
);

assign C211T=c2011T+c2111T+c2211T+c2311T+c2411T+c2511T+c2611T+c2711T+c2811T+c2911T+c2A11T+c2B11T+c2C11T+c2D11T+c2E11T+c2F11T;
assign A211T=(C211T>=0)?1:0;

assign P311T=A211T;

ninexnine_unit ninexnine_unit_7220(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2T000),
				.b1(W2T010),
				.b2(W2T020),
				.b3(W2T100),
				.b4(W2T110),
				.b5(W2T120),
				.b6(W2T200),
				.b7(W2T210),
				.b8(W2T220),
				.c(c2012T)
);

ninexnine_unit ninexnine_unit_7221(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2T001),
				.b1(W2T011),
				.b2(W2T021),
				.b3(W2T101),
				.b4(W2T111),
				.b5(W2T121),
				.b6(W2T201),
				.b7(W2T211),
				.b8(W2T221),
				.c(c2112T)
);

ninexnine_unit ninexnine_unit_7222(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2T002),
				.b1(W2T012),
				.b2(W2T022),
				.b3(W2T102),
				.b4(W2T112),
				.b5(W2T122),
				.b6(W2T202),
				.b7(W2T212),
				.b8(W2T222),
				.c(c2212T)
);

ninexnine_unit ninexnine_unit_7223(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2T003),
				.b1(W2T013),
				.b2(W2T023),
				.b3(W2T103),
				.b4(W2T113),
				.b5(W2T123),
				.b6(W2T203),
				.b7(W2T213),
				.b8(W2T223),
				.c(c2312T)
);

ninexnine_unit ninexnine_unit_7224(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2T004),
				.b1(W2T014),
				.b2(W2T024),
				.b3(W2T104),
				.b4(W2T114),
				.b5(W2T124),
				.b6(W2T204),
				.b7(W2T214),
				.b8(W2T224),
				.c(c2412T)
);

ninexnine_unit ninexnine_unit_7225(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2T005),
				.b1(W2T015),
				.b2(W2T025),
				.b3(W2T105),
				.b4(W2T115),
				.b5(W2T125),
				.b6(W2T205),
				.b7(W2T215),
				.b8(W2T225),
				.c(c2512T)
);

ninexnine_unit ninexnine_unit_7226(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2T006),
				.b1(W2T016),
				.b2(W2T026),
				.b3(W2T106),
				.b4(W2T116),
				.b5(W2T126),
				.b6(W2T206),
				.b7(W2T216),
				.b8(W2T226),
				.c(c2612T)
);

ninexnine_unit ninexnine_unit_7227(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2T007),
				.b1(W2T017),
				.b2(W2T027),
				.b3(W2T107),
				.b4(W2T117),
				.b5(W2T127),
				.b6(W2T207),
				.b7(W2T217),
				.b8(W2T227),
				.c(c2712T)
);

ninexnine_unit ninexnine_unit_7228(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2T008),
				.b1(W2T018),
				.b2(W2T028),
				.b3(W2T108),
				.b4(W2T118),
				.b5(W2T128),
				.b6(W2T208),
				.b7(W2T218),
				.b8(W2T228),
				.c(c2812T)
);

ninexnine_unit ninexnine_unit_7229(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2T009),
				.b1(W2T019),
				.b2(W2T029),
				.b3(W2T109),
				.b4(W2T119),
				.b5(W2T129),
				.b6(W2T209),
				.b7(W2T219),
				.b8(W2T229),
				.c(c2912T)
);

ninexnine_unit ninexnine_unit_7230(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2T00A),
				.b1(W2T01A),
				.b2(W2T02A),
				.b3(W2T10A),
				.b4(W2T11A),
				.b5(W2T12A),
				.b6(W2T20A),
				.b7(W2T21A),
				.b8(W2T22A),
				.c(c2A12T)
);

ninexnine_unit ninexnine_unit_7231(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2T00B),
				.b1(W2T01B),
				.b2(W2T02B),
				.b3(W2T10B),
				.b4(W2T11B),
				.b5(W2T12B),
				.b6(W2T20B),
				.b7(W2T21B),
				.b8(W2T22B),
				.c(c2B12T)
);

ninexnine_unit ninexnine_unit_7232(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2T00C),
				.b1(W2T01C),
				.b2(W2T02C),
				.b3(W2T10C),
				.b4(W2T11C),
				.b5(W2T12C),
				.b6(W2T20C),
				.b7(W2T21C),
				.b8(W2T22C),
				.c(c2C12T)
);

ninexnine_unit ninexnine_unit_7233(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2T00D),
				.b1(W2T01D),
				.b2(W2T02D),
				.b3(W2T10D),
				.b4(W2T11D),
				.b5(W2T12D),
				.b6(W2T20D),
				.b7(W2T21D),
				.b8(W2T22D),
				.c(c2D12T)
);

ninexnine_unit ninexnine_unit_7234(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2T00E),
				.b1(W2T01E),
				.b2(W2T02E),
				.b3(W2T10E),
				.b4(W2T11E),
				.b5(W2T12E),
				.b6(W2T20E),
				.b7(W2T21E),
				.b8(W2T22E),
				.c(c2E12T)
);

ninexnine_unit ninexnine_unit_7235(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2T00F),
				.b1(W2T01F),
				.b2(W2T02F),
				.b3(W2T10F),
				.b4(W2T11F),
				.b5(W2T12F),
				.b6(W2T20F),
				.b7(W2T21F),
				.b8(W2T22F),
				.c(c2F12T)
);

assign C212T=c2012T+c2112T+c2212T+c2312T+c2412T+c2512T+c2612T+c2712T+c2812T+c2912T+c2A12T+c2B12T+c2C12T+c2D12T+c2E12T+c2F12T;
assign A212T=(C212T>=0)?1:0;

assign P312T=A212T;

ninexnine_unit ninexnine_unit_7236(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2T000),
				.b1(W2T010),
				.b2(W2T020),
				.b3(W2T100),
				.b4(W2T110),
				.b5(W2T120),
				.b6(W2T200),
				.b7(W2T210),
				.b8(W2T220),
				.c(c2020T)
);

ninexnine_unit ninexnine_unit_7237(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2T001),
				.b1(W2T011),
				.b2(W2T021),
				.b3(W2T101),
				.b4(W2T111),
				.b5(W2T121),
				.b6(W2T201),
				.b7(W2T211),
				.b8(W2T221),
				.c(c2120T)
);

ninexnine_unit ninexnine_unit_7238(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2T002),
				.b1(W2T012),
				.b2(W2T022),
				.b3(W2T102),
				.b4(W2T112),
				.b5(W2T122),
				.b6(W2T202),
				.b7(W2T212),
				.b8(W2T222),
				.c(c2220T)
);

ninexnine_unit ninexnine_unit_7239(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2T003),
				.b1(W2T013),
				.b2(W2T023),
				.b3(W2T103),
				.b4(W2T113),
				.b5(W2T123),
				.b6(W2T203),
				.b7(W2T213),
				.b8(W2T223),
				.c(c2320T)
);

ninexnine_unit ninexnine_unit_7240(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2T004),
				.b1(W2T014),
				.b2(W2T024),
				.b3(W2T104),
				.b4(W2T114),
				.b5(W2T124),
				.b6(W2T204),
				.b7(W2T214),
				.b8(W2T224),
				.c(c2420T)
);

ninexnine_unit ninexnine_unit_7241(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2T005),
				.b1(W2T015),
				.b2(W2T025),
				.b3(W2T105),
				.b4(W2T115),
				.b5(W2T125),
				.b6(W2T205),
				.b7(W2T215),
				.b8(W2T225),
				.c(c2520T)
);

ninexnine_unit ninexnine_unit_7242(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2T006),
				.b1(W2T016),
				.b2(W2T026),
				.b3(W2T106),
				.b4(W2T116),
				.b5(W2T126),
				.b6(W2T206),
				.b7(W2T216),
				.b8(W2T226),
				.c(c2620T)
);

ninexnine_unit ninexnine_unit_7243(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2T007),
				.b1(W2T017),
				.b2(W2T027),
				.b3(W2T107),
				.b4(W2T117),
				.b5(W2T127),
				.b6(W2T207),
				.b7(W2T217),
				.b8(W2T227),
				.c(c2720T)
);

ninexnine_unit ninexnine_unit_7244(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2T008),
				.b1(W2T018),
				.b2(W2T028),
				.b3(W2T108),
				.b4(W2T118),
				.b5(W2T128),
				.b6(W2T208),
				.b7(W2T218),
				.b8(W2T228),
				.c(c2820T)
);

ninexnine_unit ninexnine_unit_7245(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2T009),
				.b1(W2T019),
				.b2(W2T029),
				.b3(W2T109),
				.b4(W2T119),
				.b5(W2T129),
				.b6(W2T209),
				.b7(W2T219),
				.b8(W2T229),
				.c(c2920T)
);

ninexnine_unit ninexnine_unit_7246(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2T00A),
				.b1(W2T01A),
				.b2(W2T02A),
				.b3(W2T10A),
				.b4(W2T11A),
				.b5(W2T12A),
				.b6(W2T20A),
				.b7(W2T21A),
				.b8(W2T22A),
				.c(c2A20T)
);

ninexnine_unit ninexnine_unit_7247(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2T00B),
				.b1(W2T01B),
				.b2(W2T02B),
				.b3(W2T10B),
				.b4(W2T11B),
				.b5(W2T12B),
				.b6(W2T20B),
				.b7(W2T21B),
				.b8(W2T22B),
				.c(c2B20T)
);

ninexnine_unit ninexnine_unit_7248(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2T00C),
				.b1(W2T01C),
				.b2(W2T02C),
				.b3(W2T10C),
				.b4(W2T11C),
				.b5(W2T12C),
				.b6(W2T20C),
				.b7(W2T21C),
				.b8(W2T22C),
				.c(c2C20T)
);

ninexnine_unit ninexnine_unit_7249(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2T00D),
				.b1(W2T01D),
				.b2(W2T02D),
				.b3(W2T10D),
				.b4(W2T11D),
				.b5(W2T12D),
				.b6(W2T20D),
				.b7(W2T21D),
				.b8(W2T22D),
				.c(c2D20T)
);

ninexnine_unit ninexnine_unit_7250(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2T00E),
				.b1(W2T01E),
				.b2(W2T02E),
				.b3(W2T10E),
				.b4(W2T11E),
				.b5(W2T12E),
				.b6(W2T20E),
				.b7(W2T21E),
				.b8(W2T22E),
				.c(c2E20T)
);

ninexnine_unit ninexnine_unit_7251(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2T00F),
				.b1(W2T01F),
				.b2(W2T02F),
				.b3(W2T10F),
				.b4(W2T11F),
				.b5(W2T12F),
				.b6(W2T20F),
				.b7(W2T21F),
				.b8(W2T22F),
				.c(c2F20T)
);

assign C220T=c2020T+c2120T+c2220T+c2320T+c2420T+c2520T+c2620T+c2720T+c2820T+c2920T+c2A20T+c2B20T+c2C20T+c2D20T+c2E20T+c2F20T;
assign A220T=(C220T>=0)?1:0;

assign P320T=A220T;

ninexnine_unit ninexnine_unit_7252(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2T000),
				.b1(W2T010),
				.b2(W2T020),
				.b3(W2T100),
				.b4(W2T110),
				.b5(W2T120),
				.b6(W2T200),
				.b7(W2T210),
				.b8(W2T220),
				.c(c2021T)
);

ninexnine_unit ninexnine_unit_7253(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2T001),
				.b1(W2T011),
				.b2(W2T021),
				.b3(W2T101),
				.b4(W2T111),
				.b5(W2T121),
				.b6(W2T201),
				.b7(W2T211),
				.b8(W2T221),
				.c(c2121T)
);

ninexnine_unit ninexnine_unit_7254(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2T002),
				.b1(W2T012),
				.b2(W2T022),
				.b3(W2T102),
				.b4(W2T112),
				.b5(W2T122),
				.b6(W2T202),
				.b7(W2T212),
				.b8(W2T222),
				.c(c2221T)
);

ninexnine_unit ninexnine_unit_7255(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2T003),
				.b1(W2T013),
				.b2(W2T023),
				.b3(W2T103),
				.b4(W2T113),
				.b5(W2T123),
				.b6(W2T203),
				.b7(W2T213),
				.b8(W2T223),
				.c(c2321T)
);

ninexnine_unit ninexnine_unit_7256(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2T004),
				.b1(W2T014),
				.b2(W2T024),
				.b3(W2T104),
				.b4(W2T114),
				.b5(W2T124),
				.b6(W2T204),
				.b7(W2T214),
				.b8(W2T224),
				.c(c2421T)
);

ninexnine_unit ninexnine_unit_7257(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2T005),
				.b1(W2T015),
				.b2(W2T025),
				.b3(W2T105),
				.b4(W2T115),
				.b5(W2T125),
				.b6(W2T205),
				.b7(W2T215),
				.b8(W2T225),
				.c(c2521T)
);

ninexnine_unit ninexnine_unit_7258(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2T006),
				.b1(W2T016),
				.b2(W2T026),
				.b3(W2T106),
				.b4(W2T116),
				.b5(W2T126),
				.b6(W2T206),
				.b7(W2T216),
				.b8(W2T226),
				.c(c2621T)
);

ninexnine_unit ninexnine_unit_7259(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2T007),
				.b1(W2T017),
				.b2(W2T027),
				.b3(W2T107),
				.b4(W2T117),
				.b5(W2T127),
				.b6(W2T207),
				.b7(W2T217),
				.b8(W2T227),
				.c(c2721T)
);

ninexnine_unit ninexnine_unit_7260(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2T008),
				.b1(W2T018),
				.b2(W2T028),
				.b3(W2T108),
				.b4(W2T118),
				.b5(W2T128),
				.b6(W2T208),
				.b7(W2T218),
				.b8(W2T228),
				.c(c2821T)
);

ninexnine_unit ninexnine_unit_7261(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2T009),
				.b1(W2T019),
				.b2(W2T029),
				.b3(W2T109),
				.b4(W2T119),
				.b5(W2T129),
				.b6(W2T209),
				.b7(W2T219),
				.b8(W2T229),
				.c(c2921T)
);

ninexnine_unit ninexnine_unit_7262(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2T00A),
				.b1(W2T01A),
				.b2(W2T02A),
				.b3(W2T10A),
				.b4(W2T11A),
				.b5(W2T12A),
				.b6(W2T20A),
				.b7(W2T21A),
				.b8(W2T22A),
				.c(c2A21T)
);

ninexnine_unit ninexnine_unit_7263(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2T00B),
				.b1(W2T01B),
				.b2(W2T02B),
				.b3(W2T10B),
				.b4(W2T11B),
				.b5(W2T12B),
				.b6(W2T20B),
				.b7(W2T21B),
				.b8(W2T22B),
				.c(c2B21T)
);

ninexnine_unit ninexnine_unit_7264(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2T00C),
				.b1(W2T01C),
				.b2(W2T02C),
				.b3(W2T10C),
				.b4(W2T11C),
				.b5(W2T12C),
				.b6(W2T20C),
				.b7(W2T21C),
				.b8(W2T22C),
				.c(c2C21T)
);

ninexnine_unit ninexnine_unit_7265(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2T00D),
				.b1(W2T01D),
				.b2(W2T02D),
				.b3(W2T10D),
				.b4(W2T11D),
				.b5(W2T12D),
				.b6(W2T20D),
				.b7(W2T21D),
				.b8(W2T22D),
				.c(c2D21T)
);

ninexnine_unit ninexnine_unit_7266(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2T00E),
				.b1(W2T01E),
				.b2(W2T02E),
				.b3(W2T10E),
				.b4(W2T11E),
				.b5(W2T12E),
				.b6(W2T20E),
				.b7(W2T21E),
				.b8(W2T22E),
				.c(c2E21T)
);

ninexnine_unit ninexnine_unit_7267(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2T00F),
				.b1(W2T01F),
				.b2(W2T02F),
				.b3(W2T10F),
				.b4(W2T11F),
				.b5(W2T12F),
				.b6(W2T20F),
				.b7(W2T21F),
				.b8(W2T22F),
				.c(c2F21T)
);

assign C221T=c2021T+c2121T+c2221T+c2321T+c2421T+c2521T+c2621T+c2721T+c2821T+c2921T+c2A21T+c2B21T+c2C21T+c2D21T+c2E21T+c2F21T;
assign A221T=(C221T>=0)?1:0;

assign P321T=A221T;

ninexnine_unit ninexnine_unit_7268(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2T000),
				.b1(W2T010),
				.b2(W2T020),
				.b3(W2T100),
				.b4(W2T110),
				.b5(W2T120),
				.b6(W2T200),
				.b7(W2T210),
				.b8(W2T220),
				.c(c2022T)
);

ninexnine_unit ninexnine_unit_7269(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2T001),
				.b1(W2T011),
				.b2(W2T021),
				.b3(W2T101),
				.b4(W2T111),
				.b5(W2T121),
				.b6(W2T201),
				.b7(W2T211),
				.b8(W2T221),
				.c(c2122T)
);

ninexnine_unit ninexnine_unit_7270(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2T002),
				.b1(W2T012),
				.b2(W2T022),
				.b3(W2T102),
				.b4(W2T112),
				.b5(W2T122),
				.b6(W2T202),
				.b7(W2T212),
				.b8(W2T222),
				.c(c2222T)
);

ninexnine_unit ninexnine_unit_7271(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2T003),
				.b1(W2T013),
				.b2(W2T023),
				.b3(W2T103),
				.b4(W2T113),
				.b5(W2T123),
				.b6(W2T203),
				.b7(W2T213),
				.b8(W2T223),
				.c(c2322T)
);

ninexnine_unit ninexnine_unit_7272(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2T004),
				.b1(W2T014),
				.b2(W2T024),
				.b3(W2T104),
				.b4(W2T114),
				.b5(W2T124),
				.b6(W2T204),
				.b7(W2T214),
				.b8(W2T224),
				.c(c2422T)
);

ninexnine_unit ninexnine_unit_7273(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2T005),
				.b1(W2T015),
				.b2(W2T025),
				.b3(W2T105),
				.b4(W2T115),
				.b5(W2T125),
				.b6(W2T205),
				.b7(W2T215),
				.b8(W2T225),
				.c(c2522T)
);

ninexnine_unit ninexnine_unit_7274(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2T006),
				.b1(W2T016),
				.b2(W2T026),
				.b3(W2T106),
				.b4(W2T116),
				.b5(W2T126),
				.b6(W2T206),
				.b7(W2T216),
				.b8(W2T226),
				.c(c2622T)
);

ninexnine_unit ninexnine_unit_7275(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2T007),
				.b1(W2T017),
				.b2(W2T027),
				.b3(W2T107),
				.b4(W2T117),
				.b5(W2T127),
				.b6(W2T207),
				.b7(W2T217),
				.b8(W2T227),
				.c(c2722T)
);

ninexnine_unit ninexnine_unit_7276(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2T008),
				.b1(W2T018),
				.b2(W2T028),
				.b3(W2T108),
				.b4(W2T118),
				.b5(W2T128),
				.b6(W2T208),
				.b7(W2T218),
				.b8(W2T228),
				.c(c2822T)
);

ninexnine_unit ninexnine_unit_7277(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2T009),
				.b1(W2T019),
				.b2(W2T029),
				.b3(W2T109),
				.b4(W2T119),
				.b5(W2T129),
				.b6(W2T209),
				.b7(W2T219),
				.b8(W2T229),
				.c(c2922T)
);

ninexnine_unit ninexnine_unit_7278(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2T00A),
				.b1(W2T01A),
				.b2(W2T02A),
				.b3(W2T10A),
				.b4(W2T11A),
				.b5(W2T12A),
				.b6(W2T20A),
				.b7(W2T21A),
				.b8(W2T22A),
				.c(c2A22T)
);

ninexnine_unit ninexnine_unit_7279(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2T00B),
				.b1(W2T01B),
				.b2(W2T02B),
				.b3(W2T10B),
				.b4(W2T11B),
				.b5(W2T12B),
				.b6(W2T20B),
				.b7(W2T21B),
				.b8(W2T22B),
				.c(c2B22T)
);

ninexnine_unit ninexnine_unit_7280(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2T00C),
				.b1(W2T01C),
				.b2(W2T02C),
				.b3(W2T10C),
				.b4(W2T11C),
				.b5(W2T12C),
				.b6(W2T20C),
				.b7(W2T21C),
				.b8(W2T22C),
				.c(c2C22T)
);

ninexnine_unit ninexnine_unit_7281(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2T00D),
				.b1(W2T01D),
				.b2(W2T02D),
				.b3(W2T10D),
				.b4(W2T11D),
				.b5(W2T12D),
				.b6(W2T20D),
				.b7(W2T21D),
				.b8(W2T22D),
				.c(c2D22T)
);

ninexnine_unit ninexnine_unit_7282(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2T00E),
				.b1(W2T01E),
				.b2(W2T02E),
				.b3(W2T10E),
				.b4(W2T11E),
				.b5(W2T12E),
				.b6(W2T20E),
				.b7(W2T21E),
				.b8(W2T22E),
				.c(c2E22T)
);

ninexnine_unit ninexnine_unit_7283(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2T00F),
				.b1(W2T01F),
				.b2(W2T02F),
				.b3(W2T10F),
				.b4(W2T11F),
				.b5(W2T12F),
				.b6(W2T20F),
				.b7(W2T21F),
				.b8(W2T22F),
				.c(c2F22T)
);

assign C222T=c2022T+c2122T+c2222T+c2322T+c2422T+c2522T+c2622T+c2722T+c2822T+c2922T+c2A22T+c2B22T+c2C22T+c2D22T+c2E22T+c2F22T;
assign A222T=(C222T>=0)?1:0;

assign P322T=A222T;

ninexnine_unit ninexnine_unit_7284(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2U000),
				.b1(W2U010),
				.b2(W2U020),
				.b3(W2U100),
				.b4(W2U110),
				.b5(W2U120),
				.b6(W2U200),
				.b7(W2U210),
				.b8(W2U220),
				.c(c2000U)
);

ninexnine_unit ninexnine_unit_7285(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2U001),
				.b1(W2U011),
				.b2(W2U021),
				.b3(W2U101),
				.b4(W2U111),
				.b5(W2U121),
				.b6(W2U201),
				.b7(W2U211),
				.b8(W2U221),
				.c(c2100U)
);

ninexnine_unit ninexnine_unit_7286(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2U002),
				.b1(W2U012),
				.b2(W2U022),
				.b3(W2U102),
				.b4(W2U112),
				.b5(W2U122),
				.b6(W2U202),
				.b7(W2U212),
				.b8(W2U222),
				.c(c2200U)
);

ninexnine_unit ninexnine_unit_7287(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2U003),
				.b1(W2U013),
				.b2(W2U023),
				.b3(W2U103),
				.b4(W2U113),
				.b5(W2U123),
				.b6(W2U203),
				.b7(W2U213),
				.b8(W2U223),
				.c(c2300U)
);

ninexnine_unit ninexnine_unit_7288(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2U004),
				.b1(W2U014),
				.b2(W2U024),
				.b3(W2U104),
				.b4(W2U114),
				.b5(W2U124),
				.b6(W2U204),
				.b7(W2U214),
				.b8(W2U224),
				.c(c2400U)
);

ninexnine_unit ninexnine_unit_7289(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2U005),
				.b1(W2U015),
				.b2(W2U025),
				.b3(W2U105),
				.b4(W2U115),
				.b5(W2U125),
				.b6(W2U205),
				.b7(W2U215),
				.b8(W2U225),
				.c(c2500U)
);

ninexnine_unit ninexnine_unit_7290(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2U006),
				.b1(W2U016),
				.b2(W2U026),
				.b3(W2U106),
				.b4(W2U116),
				.b5(W2U126),
				.b6(W2U206),
				.b7(W2U216),
				.b8(W2U226),
				.c(c2600U)
);

ninexnine_unit ninexnine_unit_7291(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2U007),
				.b1(W2U017),
				.b2(W2U027),
				.b3(W2U107),
				.b4(W2U117),
				.b5(W2U127),
				.b6(W2U207),
				.b7(W2U217),
				.b8(W2U227),
				.c(c2700U)
);

ninexnine_unit ninexnine_unit_7292(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2U008),
				.b1(W2U018),
				.b2(W2U028),
				.b3(W2U108),
				.b4(W2U118),
				.b5(W2U128),
				.b6(W2U208),
				.b7(W2U218),
				.b8(W2U228),
				.c(c2800U)
);

ninexnine_unit ninexnine_unit_7293(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2U009),
				.b1(W2U019),
				.b2(W2U029),
				.b3(W2U109),
				.b4(W2U119),
				.b5(W2U129),
				.b6(W2U209),
				.b7(W2U219),
				.b8(W2U229),
				.c(c2900U)
);

ninexnine_unit ninexnine_unit_7294(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2U00A),
				.b1(W2U01A),
				.b2(W2U02A),
				.b3(W2U10A),
				.b4(W2U11A),
				.b5(W2U12A),
				.b6(W2U20A),
				.b7(W2U21A),
				.b8(W2U22A),
				.c(c2A00U)
);

ninexnine_unit ninexnine_unit_7295(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2U00B),
				.b1(W2U01B),
				.b2(W2U02B),
				.b3(W2U10B),
				.b4(W2U11B),
				.b5(W2U12B),
				.b6(W2U20B),
				.b7(W2U21B),
				.b8(W2U22B),
				.c(c2B00U)
);

ninexnine_unit ninexnine_unit_7296(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2U00C),
				.b1(W2U01C),
				.b2(W2U02C),
				.b3(W2U10C),
				.b4(W2U11C),
				.b5(W2U12C),
				.b6(W2U20C),
				.b7(W2U21C),
				.b8(W2U22C),
				.c(c2C00U)
);

ninexnine_unit ninexnine_unit_7297(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2U00D),
				.b1(W2U01D),
				.b2(W2U02D),
				.b3(W2U10D),
				.b4(W2U11D),
				.b5(W2U12D),
				.b6(W2U20D),
				.b7(W2U21D),
				.b8(W2U22D),
				.c(c2D00U)
);

ninexnine_unit ninexnine_unit_7298(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2U00E),
				.b1(W2U01E),
				.b2(W2U02E),
				.b3(W2U10E),
				.b4(W2U11E),
				.b5(W2U12E),
				.b6(W2U20E),
				.b7(W2U21E),
				.b8(W2U22E),
				.c(c2E00U)
);

ninexnine_unit ninexnine_unit_7299(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2U00F),
				.b1(W2U01F),
				.b2(W2U02F),
				.b3(W2U10F),
				.b4(W2U11F),
				.b5(W2U12F),
				.b6(W2U20F),
				.b7(W2U21F),
				.b8(W2U22F),
				.c(c2F00U)
);

assign C200U=c2000U+c2100U+c2200U+c2300U+c2400U+c2500U+c2600U+c2700U+c2800U+c2900U+c2A00U+c2B00U+c2C00U+c2D00U+c2E00U+c2F00U;
assign A200U=(C200U>=0)?1:0;

assign P300U=A200U;

ninexnine_unit ninexnine_unit_7300(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2U000),
				.b1(W2U010),
				.b2(W2U020),
				.b3(W2U100),
				.b4(W2U110),
				.b5(W2U120),
				.b6(W2U200),
				.b7(W2U210),
				.b8(W2U220),
				.c(c2001U)
);

ninexnine_unit ninexnine_unit_7301(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2U001),
				.b1(W2U011),
				.b2(W2U021),
				.b3(W2U101),
				.b4(W2U111),
				.b5(W2U121),
				.b6(W2U201),
				.b7(W2U211),
				.b8(W2U221),
				.c(c2101U)
);

ninexnine_unit ninexnine_unit_7302(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2U002),
				.b1(W2U012),
				.b2(W2U022),
				.b3(W2U102),
				.b4(W2U112),
				.b5(W2U122),
				.b6(W2U202),
				.b7(W2U212),
				.b8(W2U222),
				.c(c2201U)
);

ninexnine_unit ninexnine_unit_7303(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2U003),
				.b1(W2U013),
				.b2(W2U023),
				.b3(W2U103),
				.b4(W2U113),
				.b5(W2U123),
				.b6(W2U203),
				.b7(W2U213),
				.b8(W2U223),
				.c(c2301U)
);

ninexnine_unit ninexnine_unit_7304(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2U004),
				.b1(W2U014),
				.b2(W2U024),
				.b3(W2U104),
				.b4(W2U114),
				.b5(W2U124),
				.b6(W2U204),
				.b7(W2U214),
				.b8(W2U224),
				.c(c2401U)
);

ninexnine_unit ninexnine_unit_7305(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2U005),
				.b1(W2U015),
				.b2(W2U025),
				.b3(W2U105),
				.b4(W2U115),
				.b5(W2U125),
				.b6(W2U205),
				.b7(W2U215),
				.b8(W2U225),
				.c(c2501U)
);

ninexnine_unit ninexnine_unit_7306(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2U006),
				.b1(W2U016),
				.b2(W2U026),
				.b3(W2U106),
				.b4(W2U116),
				.b5(W2U126),
				.b6(W2U206),
				.b7(W2U216),
				.b8(W2U226),
				.c(c2601U)
);

ninexnine_unit ninexnine_unit_7307(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2U007),
				.b1(W2U017),
				.b2(W2U027),
				.b3(W2U107),
				.b4(W2U117),
				.b5(W2U127),
				.b6(W2U207),
				.b7(W2U217),
				.b8(W2U227),
				.c(c2701U)
);

ninexnine_unit ninexnine_unit_7308(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2U008),
				.b1(W2U018),
				.b2(W2U028),
				.b3(W2U108),
				.b4(W2U118),
				.b5(W2U128),
				.b6(W2U208),
				.b7(W2U218),
				.b8(W2U228),
				.c(c2801U)
);

ninexnine_unit ninexnine_unit_7309(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2U009),
				.b1(W2U019),
				.b2(W2U029),
				.b3(W2U109),
				.b4(W2U119),
				.b5(W2U129),
				.b6(W2U209),
				.b7(W2U219),
				.b8(W2U229),
				.c(c2901U)
);

ninexnine_unit ninexnine_unit_7310(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2U00A),
				.b1(W2U01A),
				.b2(W2U02A),
				.b3(W2U10A),
				.b4(W2U11A),
				.b5(W2U12A),
				.b6(W2U20A),
				.b7(W2U21A),
				.b8(W2U22A),
				.c(c2A01U)
);

ninexnine_unit ninexnine_unit_7311(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2U00B),
				.b1(W2U01B),
				.b2(W2U02B),
				.b3(W2U10B),
				.b4(W2U11B),
				.b5(W2U12B),
				.b6(W2U20B),
				.b7(W2U21B),
				.b8(W2U22B),
				.c(c2B01U)
);

ninexnine_unit ninexnine_unit_7312(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2U00C),
				.b1(W2U01C),
				.b2(W2U02C),
				.b3(W2U10C),
				.b4(W2U11C),
				.b5(W2U12C),
				.b6(W2U20C),
				.b7(W2U21C),
				.b8(W2U22C),
				.c(c2C01U)
);

ninexnine_unit ninexnine_unit_7313(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2U00D),
				.b1(W2U01D),
				.b2(W2U02D),
				.b3(W2U10D),
				.b4(W2U11D),
				.b5(W2U12D),
				.b6(W2U20D),
				.b7(W2U21D),
				.b8(W2U22D),
				.c(c2D01U)
);

ninexnine_unit ninexnine_unit_7314(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2U00E),
				.b1(W2U01E),
				.b2(W2U02E),
				.b3(W2U10E),
				.b4(W2U11E),
				.b5(W2U12E),
				.b6(W2U20E),
				.b7(W2U21E),
				.b8(W2U22E),
				.c(c2E01U)
);

ninexnine_unit ninexnine_unit_7315(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2U00F),
				.b1(W2U01F),
				.b2(W2U02F),
				.b3(W2U10F),
				.b4(W2U11F),
				.b5(W2U12F),
				.b6(W2U20F),
				.b7(W2U21F),
				.b8(W2U22F),
				.c(c2F01U)
);

assign C201U=c2001U+c2101U+c2201U+c2301U+c2401U+c2501U+c2601U+c2701U+c2801U+c2901U+c2A01U+c2B01U+c2C01U+c2D01U+c2E01U+c2F01U;
assign A201U=(C201U>=0)?1:0;

assign P301U=A201U;

ninexnine_unit ninexnine_unit_7316(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2U000),
				.b1(W2U010),
				.b2(W2U020),
				.b3(W2U100),
				.b4(W2U110),
				.b5(W2U120),
				.b6(W2U200),
				.b7(W2U210),
				.b8(W2U220),
				.c(c2002U)
);

ninexnine_unit ninexnine_unit_7317(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2U001),
				.b1(W2U011),
				.b2(W2U021),
				.b3(W2U101),
				.b4(W2U111),
				.b5(W2U121),
				.b6(W2U201),
				.b7(W2U211),
				.b8(W2U221),
				.c(c2102U)
);

ninexnine_unit ninexnine_unit_7318(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2U002),
				.b1(W2U012),
				.b2(W2U022),
				.b3(W2U102),
				.b4(W2U112),
				.b5(W2U122),
				.b6(W2U202),
				.b7(W2U212),
				.b8(W2U222),
				.c(c2202U)
);

ninexnine_unit ninexnine_unit_7319(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2U003),
				.b1(W2U013),
				.b2(W2U023),
				.b3(W2U103),
				.b4(W2U113),
				.b5(W2U123),
				.b6(W2U203),
				.b7(W2U213),
				.b8(W2U223),
				.c(c2302U)
);

ninexnine_unit ninexnine_unit_7320(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2U004),
				.b1(W2U014),
				.b2(W2U024),
				.b3(W2U104),
				.b4(W2U114),
				.b5(W2U124),
				.b6(W2U204),
				.b7(W2U214),
				.b8(W2U224),
				.c(c2402U)
);

ninexnine_unit ninexnine_unit_7321(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2U005),
				.b1(W2U015),
				.b2(W2U025),
				.b3(W2U105),
				.b4(W2U115),
				.b5(W2U125),
				.b6(W2U205),
				.b7(W2U215),
				.b8(W2U225),
				.c(c2502U)
);

ninexnine_unit ninexnine_unit_7322(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2U006),
				.b1(W2U016),
				.b2(W2U026),
				.b3(W2U106),
				.b4(W2U116),
				.b5(W2U126),
				.b6(W2U206),
				.b7(W2U216),
				.b8(W2U226),
				.c(c2602U)
);

ninexnine_unit ninexnine_unit_7323(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2U007),
				.b1(W2U017),
				.b2(W2U027),
				.b3(W2U107),
				.b4(W2U117),
				.b5(W2U127),
				.b6(W2U207),
				.b7(W2U217),
				.b8(W2U227),
				.c(c2702U)
);

ninexnine_unit ninexnine_unit_7324(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2U008),
				.b1(W2U018),
				.b2(W2U028),
				.b3(W2U108),
				.b4(W2U118),
				.b5(W2U128),
				.b6(W2U208),
				.b7(W2U218),
				.b8(W2U228),
				.c(c2802U)
);

ninexnine_unit ninexnine_unit_7325(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2U009),
				.b1(W2U019),
				.b2(W2U029),
				.b3(W2U109),
				.b4(W2U119),
				.b5(W2U129),
				.b6(W2U209),
				.b7(W2U219),
				.b8(W2U229),
				.c(c2902U)
);

ninexnine_unit ninexnine_unit_7326(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2U00A),
				.b1(W2U01A),
				.b2(W2U02A),
				.b3(W2U10A),
				.b4(W2U11A),
				.b5(W2U12A),
				.b6(W2U20A),
				.b7(W2U21A),
				.b8(W2U22A),
				.c(c2A02U)
);

ninexnine_unit ninexnine_unit_7327(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2U00B),
				.b1(W2U01B),
				.b2(W2U02B),
				.b3(W2U10B),
				.b4(W2U11B),
				.b5(W2U12B),
				.b6(W2U20B),
				.b7(W2U21B),
				.b8(W2U22B),
				.c(c2B02U)
);

ninexnine_unit ninexnine_unit_7328(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2U00C),
				.b1(W2U01C),
				.b2(W2U02C),
				.b3(W2U10C),
				.b4(W2U11C),
				.b5(W2U12C),
				.b6(W2U20C),
				.b7(W2U21C),
				.b8(W2U22C),
				.c(c2C02U)
);

ninexnine_unit ninexnine_unit_7329(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2U00D),
				.b1(W2U01D),
				.b2(W2U02D),
				.b3(W2U10D),
				.b4(W2U11D),
				.b5(W2U12D),
				.b6(W2U20D),
				.b7(W2U21D),
				.b8(W2U22D),
				.c(c2D02U)
);

ninexnine_unit ninexnine_unit_7330(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2U00E),
				.b1(W2U01E),
				.b2(W2U02E),
				.b3(W2U10E),
				.b4(W2U11E),
				.b5(W2U12E),
				.b6(W2U20E),
				.b7(W2U21E),
				.b8(W2U22E),
				.c(c2E02U)
);

ninexnine_unit ninexnine_unit_7331(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2U00F),
				.b1(W2U01F),
				.b2(W2U02F),
				.b3(W2U10F),
				.b4(W2U11F),
				.b5(W2U12F),
				.b6(W2U20F),
				.b7(W2U21F),
				.b8(W2U22F),
				.c(c2F02U)
);

assign C202U=c2002U+c2102U+c2202U+c2302U+c2402U+c2502U+c2602U+c2702U+c2802U+c2902U+c2A02U+c2B02U+c2C02U+c2D02U+c2E02U+c2F02U;
assign A202U=(C202U>=0)?1:0;

assign P302U=A202U;

ninexnine_unit ninexnine_unit_7332(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2U000),
				.b1(W2U010),
				.b2(W2U020),
				.b3(W2U100),
				.b4(W2U110),
				.b5(W2U120),
				.b6(W2U200),
				.b7(W2U210),
				.b8(W2U220),
				.c(c2010U)
);

ninexnine_unit ninexnine_unit_7333(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2U001),
				.b1(W2U011),
				.b2(W2U021),
				.b3(W2U101),
				.b4(W2U111),
				.b5(W2U121),
				.b6(W2U201),
				.b7(W2U211),
				.b8(W2U221),
				.c(c2110U)
);

ninexnine_unit ninexnine_unit_7334(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2U002),
				.b1(W2U012),
				.b2(W2U022),
				.b3(W2U102),
				.b4(W2U112),
				.b5(W2U122),
				.b6(W2U202),
				.b7(W2U212),
				.b8(W2U222),
				.c(c2210U)
);

ninexnine_unit ninexnine_unit_7335(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2U003),
				.b1(W2U013),
				.b2(W2U023),
				.b3(W2U103),
				.b4(W2U113),
				.b5(W2U123),
				.b6(W2U203),
				.b7(W2U213),
				.b8(W2U223),
				.c(c2310U)
);

ninexnine_unit ninexnine_unit_7336(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2U004),
				.b1(W2U014),
				.b2(W2U024),
				.b3(W2U104),
				.b4(W2U114),
				.b5(W2U124),
				.b6(W2U204),
				.b7(W2U214),
				.b8(W2U224),
				.c(c2410U)
);

ninexnine_unit ninexnine_unit_7337(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2U005),
				.b1(W2U015),
				.b2(W2U025),
				.b3(W2U105),
				.b4(W2U115),
				.b5(W2U125),
				.b6(W2U205),
				.b7(W2U215),
				.b8(W2U225),
				.c(c2510U)
);

ninexnine_unit ninexnine_unit_7338(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2U006),
				.b1(W2U016),
				.b2(W2U026),
				.b3(W2U106),
				.b4(W2U116),
				.b5(W2U126),
				.b6(W2U206),
				.b7(W2U216),
				.b8(W2U226),
				.c(c2610U)
);

ninexnine_unit ninexnine_unit_7339(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2U007),
				.b1(W2U017),
				.b2(W2U027),
				.b3(W2U107),
				.b4(W2U117),
				.b5(W2U127),
				.b6(W2U207),
				.b7(W2U217),
				.b8(W2U227),
				.c(c2710U)
);

ninexnine_unit ninexnine_unit_7340(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2U008),
				.b1(W2U018),
				.b2(W2U028),
				.b3(W2U108),
				.b4(W2U118),
				.b5(W2U128),
				.b6(W2U208),
				.b7(W2U218),
				.b8(W2U228),
				.c(c2810U)
);

ninexnine_unit ninexnine_unit_7341(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2U009),
				.b1(W2U019),
				.b2(W2U029),
				.b3(W2U109),
				.b4(W2U119),
				.b5(W2U129),
				.b6(W2U209),
				.b7(W2U219),
				.b8(W2U229),
				.c(c2910U)
);

ninexnine_unit ninexnine_unit_7342(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2U00A),
				.b1(W2U01A),
				.b2(W2U02A),
				.b3(W2U10A),
				.b4(W2U11A),
				.b5(W2U12A),
				.b6(W2U20A),
				.b7(W2U21A),
				.b8(W2U22A),
				.c(c2A10U)
);

ninexnine_unit ninexnine_unit_7343(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2U00B),
				.b1(W2U01B),
				.b2(W2U02B),
				.b3(W2U10B),
				.b4(W2U11B),
				.b5(W2U12B),
				.b6(W2U20B),
				.b7(W2U21B),
				.b8(W2U22B),
				.c(c2B10U)
);

ninexnine_unit ninexnine_unit_7344(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2U00C),
				.b1(W2U01C),
				.b2(W2U02C),
				.b3(W2U10C),
				.b4(W2U11C),
				.b5(W2U12C),
				.b6(W2U20C),
				.b7(W2U21C),
				.b8(W2U22C),
				.c(c2C10U)
);

ninexnine_unit ninexnine_unit_7345(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2U00D),
				.b1(W2U01D),
				.b2(W2U02D),
				.b3(W2U10D),
				.b4(W2U11D),
				.b5(W2U12D),
				.b6(W2U20D),
				.b7(W2U21D),
				.b8(W2U22D),
				.c(c2D10U)
);

ninexnine_unit ninexnine_unit_7346(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2U00E),
				.b1(W2U01E),
				.b2(W2U02E),
				.b3(W2U10E),
				.b4(W2U11E),
				.b5(W2U12E),
				.b6(W2U20E),
				.b7(W2U21E),
				.b8(W2U22E),
				.c(c2E10U)
);

ninexnine_unit ninexnine_unit_7347(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2U00F),
				.b1(W2U01F),
				.b2(W2U02F),
				.b3(W2U10F),
				.b4(W2U11F),
				.b5(W2U12F),
				.b6(W2U20F),
				.b7(W2U21F),
				.b8(W2U22F),
				.c(c2F10U)
);

assign C210U=c2010U+c2110U+c2210U+c2310U+c2410U+c2510U+c2610U+c2710U+c2810U+c2910U+c2A10U+c2B10U+c2C10U+c2D10U+c2E10U+c2F10U;
assign A210U=(C210U>=0)?1:0;

assign P310U=A210U;

ninexnine_unit ninexnine_unit_7348(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2U000),
				.b1(W2U010),
				.b2(W2U020),
				.b3(W2U100),
				.b4(W2U110),
				.b5(W2U120),
				.b6(W2U200),
				.b7(W2U210),
				.b8(W2U220),
				.c(c2011U)
);

ninexnine_unit ninexnine_unit_7349(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2U001),
				.b1(W2U011),
				.b2(W2U021),
				.b3(W2U101),
				.b4(W2U111),
				.b5(W2U121),
				.b6(W2U201),
				.b7(W2U211),
				.b8(W2U221),
				.c(c2111U)
);

ninexnine_unit ninexnine_unit_7350(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2U002),
				.b1(W2U012),
				.b2(W2U022),
				.b3(W2U102),
				.b4(W2U112),
				.b5(W2U122),
				.b6(W2U202),
				.b7(W2U212),
				.b8(W2U222),
				.c(c2211U)
);

ninexnine_unit ninexnine_unit_7351(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2U003),
				.b1(W2U013),
				.b2(W2U023),
				.b3(W2U103),
				.b4(W2U113),
				.b5(W2U123),
				.b6(W2U203),
				.b7(W2U213),
				.b8(W2U223),
				.c(c2311U)
);

ninexnine_unit ninexnine_unit_7352(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2U004),
				.b1(W2U014),
				.b2(W2U024),
				.b3(W2U104),
				.b4(W2U114),
				.b5(W2U124),
				.b6(W2U204),
				.b7(W2U214),
				.b8(W2U224),
				.c(c2411U)
);

ninexnine_unit ninexnine_unit_7353(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2U005),
				.b1(W2U015),
				.b2(W2U025),
				.b3(W2U105),
				.b4(W2U115),
				.b5(W2U125),
				.b6(W2U205),
				.b7(W2U215),
				.b8(W2U225),
				.c(c2511U)
);

ninexnine_unit ninexnine_unit_7354(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2U006),
				.b1(W2U016),
				.b2(W2U026),
				.b3(W2U106),
				.b4(W2U116),
				.b5(W2U126),
				.b6(W2U206),
				.b7(W2U216),
				.b8(W2U226),
				.c(c2611U)
);

ninexnine_unit ninexnine_unit_7355(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2U007),
				.b1(W2U017),
				.b2(W2U027),
				.b3(W2U107),
				.b4(W2U117),
				.b5(W2U127),
				.b6(W2U207),
				.b7(W2U217),
				.b8(W2U227),
				.c(c2711U)
);

ninexnine_unit ninexnine_unit_7356(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2U008),
				.b1(W2U018),
				.b2(W2U028),
				.b3(W2U108),
				.b4(W2U118),
				.b5(W2U128),
				.b6(W2U208),
				.b7(W2U218),
				.b8(W2U228),
				.c(c2811U)
);

ninexnine_unit ninexnine_unit_7357(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2U009),
				.b1(W2U019),
				.b2(W2U029),
				.b3(W2U109),
				.b4(W2U119),
				.b5(W2U129),
				.b6(W2U209),
				.b7(W2U219),
				.b8(W2U229),
				.c(c2911U)
);

ninexnine_unit ninexnine_unit_7358(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2U00A),
				.b1(W2U01A),
				.b2(W2U02A),
				.b3(W2U10A),
				.b4(W2U11A),
				.b5(W2U12A),
				.b6(W2U20A),
				.b7(W2U21A),
				.b8(W2U22A),
				.c(c2A11U)
);

ninexnine_unit ninexnine_unit_7359(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2U00B),
				.b1(W2U01B),
				.b2(W2U02B),
				.b3(W2U10B),
				.b4(W2U11B),
				.b5(W2U12B),
				.b6(W2U20B),
				.b7(W2U21B),
				.b8(W2U22B),
				.c(c2B11U)
);

ninexnine_unit ninexnine_unit_7360(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2U00C),
				.b1(W2U01C),
				.b2(W2U02C),
				.b3(W2U10C),
				.b4(W2U11C),
				.b5(W2U12C),
				.b6(W2U20C),
				.b7(W2U21C),
				.b8(W2U22C),
				.c(c2C11U)
);

ninexnine_unit ninexnine_unit_7361(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2U00D),
				.b1(W2U01D),
				.b2(W2U02D),
				.b3(W2U10D),
				.b4(W2U11D),
				.b5(W2U12D),
				.b6(W2U20D),
				.b7(W2U21D),
				.b8(W2U22D),
				.c(c2D11U)
);

ninexnine_unit ninexnine_unit_7362(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2U00E),
				.b1(W2U01E),
				.b2(W2U02E),
				.b3(W2U10E),
				.b4(W2U11E),
				.b5(W2U12E),
				.b6(W2U20E),
				.b7(W2U21E),
				.b8(W2U22E),
				.c(c2E11U)
);

ninexnine_unit ninexnine_unit_7363(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2U00F),
				.b1(W2U01F),
				.b2(W2U02F),
				.b3(W2U10F),
				.b4(W2U11F),
				.b5(W2U12F),
				.b6(W2U20F),
				.b7(W2U21F),
				.b8(W2U22F),
				.c(c2F11U)
);

assign C211U=c2011U+c2111U+c2211U+c2311U+c2411U+c2511U+c2611U+c2711U+c2811U+c2911U+c2A11U+c2B11U+c2C11U+c2D11U+c2E11U+c2F11U;
assign A211U=(C211U>=0)?1:0;

assign P311U=A211U;

ninexnine_unit ninexnine_unit_7364(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2U000),
				.b1(W2U010),
				.b2(W2U020),
				.b3(W2U100),
				.b4(W2U110),
				.b5(W2U120),
				.b6(W2U200),
				.b7(W2U210),
				.b8(W2U220),
				.c(c2012U)
);

ninexnine_unit ninexnine_unit_7365(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2U001),
				.b1(W2U011),
				.b2(W2U021),
				.b3(W2U101),
				.b4(W2U111),
				.b5(W2U121),
				.b6(W2U201),
				.b7(W2U211),
				.b8(W2U221),
				.c(c2112U)
);

ninexnine_unit ninexnine_unit_7366(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2U002),
				.b1(W2U012),
				.b2(W2U022),
				.b3(W2U102),
				.b4(W2U112),
				.b5(W2U122),
				.b6(W2U202),
				.b7(W2U212),
				.b8(W2U222),
				.c(c2212U)
);

ninexnine_unit ninexnine_unit_7367(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2U003),
				.b1(W2U013),
				.b2(W2U023),
				.b3(W2U103),
				.b4(W2U113),
				.b5(W2U123),
				.b6(W2U203),
				.b7(W2U213),
				.b8(W2U223),
				.c(c2312U)
);

ninexnine_unit ninexnine_unit_7368(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2U004),
				.b1(W2U014),
				.b2(W2U024),
				.b3(W2U104),
				.b4(W2U114),
				.b5(W2U124),
				.b6(W2U204),
				.b7(W2U214),
				.b8(W2U224),
				.c(c2412U)
);

ninexnine_unit ninexnine_unit_7369(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2U005),
				.b1(W2U015),
				.b2(W2U025),
				.b3(W2U105),
				.b4(W2U115),
				.b5(W2U125),
				.b6(W2U205),
				.b7(W2U215),
				.b8(W2U225),
				.c(c2512U)
);

ninexnine_unit ninexnine_unit_7370(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2U006),
				.b1(W2U016),
				.b2(W2U026),
				.b3(W2U106),
				.b4(W2U116),
				.b5(W2U126),
				.b6(W2U206),
				.b7(W2U216),
				.b8(W2U226),
				.c(c2612U)
);

ninexnine_unit ninexnine_unit_7371(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2U007),
				.b1(W2U017),
				.b2(W2U027),
				.b3(W2U107),
				.b4(W2U117),
				.b5(W2U127),
				.b6(W2U207),
				.b7(W2U217),
				.b8(W2U227),
				.c(c2712U)
);

ninexnine_unit ninexnine_unit_7372(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2U008),
				.b1(W2U018),
				.b2(W2U028),
				.b3(W2U108),
				.b4(W2U118),
				.b5(W2U128),
				.b6(W2U208),
				.b7(W2U218),
				.b8(W2U228),
				.c(c2812U)
);

ninexnine_unit ninexnine_unit_7373(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2U009),
				.b1(W2U019),
				.b2(W2U029),
				.b3(W2U109),
				.b4(W2U119),
				.b5(W2U129),
				.b6(W2U209),
				.b7(W2U219),
				.b8(W2U229),
				.c(c2912U)
);

ninexnine_unit ninexnine_unit_7374(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2U00A),
				.b1(W2U01A),
				.b2(W2U02A),
				.b3(W2U10A),
				.b4(W2U11A),
				.b5(W2U12A),
				.b6(W2U20A),
				.b7(W2U21A),
				.b8(W2U22A),
				.c(c2A12U)
);

ninexnine_unit ninexnine_unit_7375(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2U00B),
				.b1(W2U01B),
				.b2(W2U02B),
				.b3(W2U10B),
				.b4(W2U11B),
				.b5(W2U12B),
				.b6(W2U20B),
				.b7(W2U21B),
				.b8(W2U22B),
				.c(c2B12U)
);

ninexnine_unit ninexnine_unit_7376(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2U00C),
				.b1(W2U01C),
				.b2(W2U02C),
				.b3(W2U10C),
				.b4(W2U11C),
				.b5(W2U12C),
				.b6(W2U20C),
				.b7(W2U21C),
				.b8(W2U22C),
				.c(c2C12U)
);

ninexnine_unit ninexnine_unit_7377(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2U00D),
				.b1(W2U01D),
				.b2(W2U02D),
				.b3(W2U10D),
				.b4(W2U11D),
				.b5(W2U12D),
				.b6(W2U20D),
				.b7(W2U21D),
				.b8(W2U22D),
				.c(c2D12U)
);

ninexnine_unit ninexnine_unit_7378(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2U00E),
				.b1(W2U01E),
				.b2(W2U02E),
				.b3(W2U10E),
				.b4(W2U11E),
				.b5(W2U12E),
				.b6(W2U20E),
				.b7(W2U21E),
				.b8(W2U22E),
				.c(c2E12U)
);

ninexnine_unit ninexnine_unit_7379(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2U00F),
				.b1(W2U01F),
				.b2(W2U02F),
				.b3(W2U10F),
				.b4(W2U11F),
				.b5(W2U12F),
				.b6(W2U20F),
				.b7(W2U21F),
				.b8(W2U22F),
				.c(c2F12U)
);

assign C212U=c2012U+c2112U+c2212U+c2312U+c2412U+c2512U+c2612U+c2712U+c2812U+c2912U+c2A12U+c2B12U+c2C12U+c2D12U+c2E12U+c2F12U;
assign A212U=(C212U>=0)?1:0;

assign P312U=A212U;

ninexnine_unit ninexnine_unit_7380(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2U000),
				.b1(W2U010),
				.b2(W2U020),
				.b3(W2U100),
				.b4(W2U110),
				.b5(W2U120),
				.b6(W2U200),
				.b7(W2U210),
				.b8(W2U220),
				.c(c2020U)
);

ninexnine_unit ninexnine_unit_7381(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2U001),
				.b1(W2U011),
				.b2(W2U021),
				.b3(W2U101),
				.b4(W2U111),
				.b5(W2U121),
				.b6(W2U201),
				.b7(W2U211),
				.b8(W2U221),
				.c(c2120U)
);

ninexnine_unit ninexnine_unit_7382(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2U002),
				.b1(W2U012),
				.b2(W2U022),
				.b3(W2U102),
				.b4(W2U112),
				.b5(W2U122),
				.b6(W2U202),
				.b7(W2U212),
				.b8(W2U222),
				.c(c2220U)
);

ninexnine_unit ninexnine_unit_7383(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2U003),
				.b1(W2U013),
				.b2(W2U023),
				.b3(W2U103),
				.b4(W2U113),
				.b5(W2U123),
				.b6(W2U203),
				.b7(W2U213),
				.b8(W2U223),
				.c(c2320U)
);

ninexnine_unit ninexnine_unit_7384(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2U004),
				.b1(W2U014),
				.b2(W2U024),
				.b3(W2U104),
				.b4(W2U114),
				.b5(W2U124),
				.b6(W2U204),
				.b7(W2U214),
				.b8(W2U224),
				.c(c2420U)
);

ninexnine_unit ninexnine_unit_7385(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2U005),
				.b1(W2U015),
				.b2(W2U025),
				.b3(W2U105),
				.b4(W2U115),
				.b5(W2U125),
				.b6(W2U205),
				.b7(W2U215),
				.b8(W2U225),
				.c(c2520U)
);

ninexnine_unit ninexnine_unit_7386(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2U006),
				.b1(W2U016),
				.b2(W2U026),
				.b3(W2U106),
				.b4(W2U116),
				.b5(W2U126),
				.b6(W2U206),
				.b7(W2U216),
				.b8(W2U226),
				.c(c2620U)
);

ninexnine_unit ninexnine_unit_7387(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2U007),
				.b1(W2U017),
				.b2(W2U027),
				.b3(W2U107),
				.b4(W2U117),
				.b5(W2U127),
				.b6(W2U207),
				.b7(W2U217),
				.b8(W2U227),
				.c(c2720U)
);

ninexnine_unit ninexnine_unit_7388(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2U008),
				.b1(W2U018),
				.b2(W2U028),
				.b3(W2U108),
				.b4(W2U118),
				.b5(W2U128),
				.b6(W2U208),
				.b7(W2U218),
				.b8(W2U228),
				.c(c2820U)
);

ninexnine_unit ninexnine_unit_7389(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2U009),
				.b1(W2U019),
				.b2(W2U029),
				.b3(W2U109),
				.b4(W2U119),
				.b5(W2U129),
				.b6(W2U209),
				.b7(W2U219),
				.b8(W2U229),
				.c(c2920U)
);

ninexnine_unit ninexnine_unit_7390(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2U00A),
				.b1(W2U01A),
				.b2(W2U02A),
				.b3(W2U10A),
				.b4(W2U11A),
				.b5(W2U12A),
				.b6(W2U20A),
				.b7(W2U21A),
				.b8(W2U22A),
				.c(c2A20U)
);

ninexnine_unit ninexnine_unit_7391(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2U00B),
				.b1(W2U01B),
				.b2(W2U02B),
				.b3(W2U10B),
				.b4(W2U11B),
				.b5(W2U12B),
				.b6(W2U20B),
				.b7(W2U21B),
				.b8(W2U22B),
				.c(c2B20U)
);

ninexnine_unit ninexnine_unit_7392(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2U00C),
				.b1(W2U01C),
				.b2(W2U02C),
				.b3(W2U10C),
				.b4(W2U11C),
				.b5(W2U12C),
				.b6(W2U20C),
				.b7(W2U21C),
				.b8(W2U22C),
				.c(c2C20U)
);

ninexnine_unit ninexnine_unit_7393(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2U00D),
				.b1(W2U01D),
				.b2(W2U02D),
				.b3(W2U10D),
				.b4(W2U11D),
				.b5(W2U12D),
				.b6(W2U20D),
				.b7(W2U21D),
				.b8(W2U22D),
				.c(c2D20U)
);

ninexnine_unit ninexnine_unit_7394(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2U00E),
				.b1(W2U01E),
				.b2(W2U02E),
				.b3(W2U10E),
				.b4(W2U11E),
				.b5(W2U12E),
				.b6(W2U20E),
				.b7(W2U21E),
				.b8(W2U22E),
				.c(c2E20U)
);

ninexnine_unit ninexnine_unit_7395(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2U00F),
				.b1(W2U01F),
				.b2(W2U02F),
				.b3(W2U10F),
				.b4(W2U11F),
				.b5(W2U12F),
				.b6(W2U20F),
				.b7(W2U21F),
				.b8(W2U22F),
				.c(c2F20U)
);

assign C220U=c2020U+c2120U+c2220U+c2320U+c2420U+c2520U+c2620U+c2720U+c2820U+c2920U+c2A20U+c2B20U+c2C20U+c2D20U+c2E20U+c2F20U;
assign A220U=(C220U>=0)?1:0;

assign P320U=A220U;

ninexnine_unit ninexnine_unit_7396(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2U000),
				.b1(W2U010),
				.b2(W2U020),
				.b3(W2U100),
				.b4(W2U110),
				.b5(W2U120),
				.b6(W2U200),
				.b7(W2U210),
				.b8(W2U220),
				.c(c2021U)
);

ninexnine_unit ninexnine_unit_7397(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2U001),
				.b1(W2U011),
				.b2(W2U021),
				.b3(W2U101),
				.b4(W2U111),
				.b5(W2U121),
				.b6(W2U201),
				.b7(W2U211),
				.b8(W2U221),
				.c(c2121U)
);

ninexnine_unit ninexnine_unit_7398(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2U002),
				.b1(W2U012),
				.b2(W2U022),
				.b3(W2U102),
				.b4(W2U112),
				.b5(W2U122),
				.b6(W2U202),
				.b7(W2U212),
				.b8(W2U222),
				.c(c2221U)
);

ninexnine_unit ninexnine_unit_7399(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2U003),
				.b1(W2U013),
				.b2(W2U023),
				.b3(W2U103),
				.b4(W2U113),
				.b5(W2U123),
				.b6(W2U203),
				.b7(W2U213),
				.b8(W2U223),
				.c(c2321U)
);

ninexnine_unit ninexnine_unit_7400(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2U004),
				.b1(W2U014),
				.b2(W2U024),
				.b3(W2U104),
				.b4(W2U114),
				.b5(W2U124),
				.b6(W2U204),
				.b7(W2U214),
				.b8(W2U224),
				.c(c2421U)
);

ninexnine_unit ninexnine_unit_7401(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2U005),
				.b1(W2U015),
				.b2(W2U025),
				.b3(W2U105),
				.b4(W2U115),
				.b5(W2U125),
				.b6(W2U205),
				.b7(W2U215),
				.b8(W2U225),
				.c(c2521U)
);

ninexnine_unit ninexnine_unit_7402(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2U006),
				.b1(W2U016),
				.b2(W2U026),
				.b3(W2U106),
				.b4(W2U116),
				.b5(W2U126),
				.b6(W2U206),
				.b7(W2U216),
				.b8(W2U226),
				.c(c2621U)
);

ninexnine_unit ninexnine_unit_7403(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2U007),
				.b1(W2U017),
				.b2(W2U027),
				.b3(W2U107),
				.b4(W2U117),
				.b5(W2U127),
				.b6(W2U207),
				.b7(W2U217),
				.b8(W2U227),
				.c(c2721U)
);

ninexnine_unit ninexnine_unit_7404(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2U008),
				.b1(W2U018),
				.b2(W2U028),
				.b3(W2U108),
				.b4(W2U118),
				.b5(W2U128),
				.b6(W2U208),
				.b7(W2U218),
				.b8(W2U228),
				.c(c2821U)
);

ninexnine_unit ninexnine_unit_7405(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2U009),
				.b1(W2U019),
				.b2(W2U029),
				.b3(W2U109),
				.b4(W2U119),
				.b5(W2U129),
				.b6(W2U209),
				.b7(W2U219),
				.b8(W2U229),
				.c(c2921U)
);

ninexnine_unit ninexnine_unit_7406(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2U00A),
				.b1(W2U01A),
				.b2(W2U02A),
				.b3(W2U10A),
				.b4(W2U11A),
				.b5(W2U12A),
				.b6(W2U20A),
				.b7(W2U21A),
				.b8(W2U22A),
				.c(c2A21U)
);

ninexnine_unit ninexnine_unit_7407(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2U00B),
				.b1(W2U01B),
				.b2(W2U02B),
				.b3(W2U10B),
				.b4(W2U11B),
				.b5(W2U12B),
				.b6(W2U20B),
				.b7(W2U21B),
				.b8(W2U22B),
				.c(c2B21U)
);

ninexnine_unit ninexnine_unit_7408(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2U00C),
				.b1(W2U01C),
				.b2(W2U02C),
				.b3(W2U10C),
				.b4(W2U11C),
				.b5(W2U12C),
				.b6(W2U20C),
				.b7(W2U21C),
				.b8(W2U22C),
				.c(c2C21U)
);

ninexnine_unit ninexnine_unit_7409(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2U00D),
				.b1(W2U01D),
				.b2(W2U02D),
				.b3(W2U10D),
				.b4(W2U11D),
				.b5(W2U12D),
				.b6(W2U20D),
				.b7(W2U21D),
				.b8(W2U22D),
				.c(c2D21U)
);

ninexnine_unit ninexnine_unit_7410(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2U00E),
				.b1(W2U01E),
				.b2(W2U02E),
				.b3(W2U10E),
				.b4(W2U11E),
				.b5(W2U12E),
				.b6(W2U20E),
				.b7(W2U21E),
				.b8(W2U22E),
				.c(c2E21U)
);

ninexnine_unit ninexnine_unit_7411(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2U00F),
				.b1(W2U01F),
				.b2(W2U02F),
				.b3(W2U10F),
				.b4(W2U11F),
				.b5(W2U12F),
				.b6(W2U20F),
				.b7(W2U21F),
				.b8(W2U22F),
				.c(c2F21U)
);

assign C221U=c2021U+c2121U+c2221U+c2321U+c2421U+c2521U+c2621U+c2721U+c2821U+c2921U+c2A21U+c2B21U+c2C21U+c2D21U+c2E21U+c2F21U;
assign A221U=(C221U>=0)?1:0;

assign P321U=A221U;

ninexnine_unit ninexnine_unit_7412(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2U000),
				.b1(W2U010),
				.b2(W2U020),
				.b3(W2U100),
				.b4(W2U110),
				.b5(W2U120),
				.b6(W2U200),
				.b7(W2U210),
				.b8(W2U220),
				.c(c2022U)
);

ninexnine_unit ninexnine_unit_7413(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2U001),
				.b1(W2U011),
				.b2(W2U021),
				.b3(W2U101),
				.b4(W2U111),
				.b5(W2U121),
				.b6(W2U201),
				.b7(W2U211),
				.b8(W2U221),
				.c(c2122U)
);

ninexnine_unit ninexnine_unit_7414(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2U002),
				.b1(W2U012),
				.b2(W2U022),
				.b3(W2U102),
				.b4(W2U112),
				.b5(W2U122),
				.b6(W2U202),
				.b7(W2U212),
				.b8(W2U222),
				.c(c2222U)
);

ninexnine_unit ninexnine_unit_7415(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2U003),
				.b1(W2U013),
				.b2(W2U023),
				.b3(W2U103),
				.b4(W2U113),
				.b5(W2U123),
				.b6(W2U203),
				.b7(W2U213),
				.b8(W2U223),
				.c(c2322U)
);

ninexnine_unit ninexnine_unit_7416(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2U004),
				.b1(W2U014),
				.b2(W2U024),
				.b3(W2U104),
				.b4(W2U114),
				.b5(W2U124),
				.b6(W2U204),
				.b7(W2U214),
				.b8(W2U224),
				.c(c2422U)
);

ninexnine_unit ninexnine_unit_7417(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2U005),
				.b1(W2U015),
				.b2(W2U025),
				.b3(W2U105),
				.b4(W2U115),
				.b5(W2U125),
				.b6(W2U205),
				.b7(W2U215),
				.b8(W2U225),
				.c(c2522U)
);

ninexnine_unit ninexnine_unit_7418(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2U006),
				.b1(W2U016),
				.b2(W2U026),
				.b3(W2U106),
				.b4(W2U116),
				.b5(W2U126),
				.b6(W2U206),
				.b7(W2U216),
				.b8(W2U226),
				.c(c2622U)
);

ninexnine_unit ninexnine_unit_7419(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2U007),
				.b1(W2U017),
				.b2(W2U027),
				.b3(W2U107),
				.b4(W2U117),
				.b5(W2U127),
				.b6(W2U207),
				.b7(W2U217),
				.b8(W2U227),
				.c(c2722U)
);

ninexnine_unit ninexnine_unit_7420(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2U008),
				.b1(W2U018),
				.b2(W2U028),
				.b3(W2U108),
				.b4(W2U118),
				.b5(W2U128),
				.b6(W2U208),
				.b7(W2U218),
				.b8(W2U228),
				.c(c2822U)
);

ninexnine_unit ninexnine_unit_7421(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2U009),
				.b1(W2U019),
				.b2(W2U029),
				.b3(W2U109),
				.b4(W2U119),
				.b5(W2U129),
				.b6(W2U209),
				.b7(W2U219),
				.b8(W2U229),
				.c(c2922U)
);

ninexnine_unit ninexnine_unit_7422(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2U00A),
				.b1(W2U01A),
				.b2(W2U02A),
				.b3(W2U10A),
				.b4(W2U11A),
				.b5(W2U12A),
				.b6(W2U20A),
				.b7(W2U21A),
				.b8(W2U22A),
				.c(c2A22U)
);

ninexnine_unit ninexnine_unit_7423(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2U00B),
				.b1(W2U01B),
				.b2(W2U02B),
				.b3(W2U10B),
				.b4(W2U11B),
				.b5(W2U12B),
				.b6(W2U20B),
				.b7(W2U21B),
				.b8(W2U22B),
				.c(c2B22U)
);

ninexnine_unit ninexnine_unit_7424(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2U00C),
				.b1(W2U01C),
				.b2(W2U02C),
				.b3(W2U10C),
				.b4(W2U11C),
				.b5(W2U12C),
				.b6(W2U20C),
				.b7(W2U21C),
				.b8(W2U22C),
				.c(c2C22U)
);

ninexnine_unit ninexnine_unit_7425(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2U00D),
				.b1(W2U01D),
				.b2(W2U02D),
				.b3(W2U10D),
				.b4(W2U11D),
				.b5(W2U12D),
				.b6(W2U20D),
				.b7(W2U21D),
				.b8(W2U22D),
				.c(c2D22U)
);

ninexnine_unit ninexnine_unit_7426(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2U00E),
				.b1(W2U01E),
				.b2(W2U02E),
				.b3(W2U10E),
				.b4(W2U11E),
				.b5(W2U12E),
				.b6(W2U20E),
				.b7(W2U21E),
				.b8(W2U22E),
				.c(c2E22U)
);

ninexnine_unit ninexnine_unit_7427(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2U00F),
				.b1(W2U01F),
				.b2(W2U02F),
				.b3(W2U10F),
				.b4(W2U11F),
				.b5(W2U12F),
				.b6(W2U20F),
				.b7(W2U21F),
				.b8(W2U22F),
				.c(c2F22U)
);

assign C222U=c2022U+c2122U+c2222U+c2322U+c2422U+c2522U+c2622U+c2722U+c2822U+c2922U+c2A22U+c2B22U+c2C22U+c2D22U+c2E22U+c2F22U;
assign A222U=(C222U>=0)?1:0;

assign P322U=A222U;

ninexnine_unit ninexnine_unit_7428(
				.clk(clk),
				.rstn(rstn),
				.a0(P2000),
				.a1(P2010),
				.a2(P2020),
				.a3(P2100),
				.a4(P2110),
				.a5(P2120),
				.a6(P2200),
				.a7(P2210),
				.a8(P2220),
				.b0(W2V000),
				.b1(W2V010),
				.b2(W2V020),
				.b3(W2V100),
				.b4(W2V110),
				.b5(W2V120),
				.b6(W2V200),
				.b7(W2V210),
				.b8(W2V220),
				.c(c2000V)
);

ninexnine_unit ninexnine_unit_7429(
				.clk(clk),
				.rstn(rstn),
				.a0(P2001),
				.a1(P2011),
				.a2(P2021),
				.a3(P2101),
				.a4(P2111),
				.a5(P2121),
				.a6(P2201),
				.a7(P2211),
				.a8(P2221),
				.b0(W2V001),
				.b1(W2V011),
				.b2(W2V021),
				.b3(W2V101),
				.b4(W2V111),
				.b5(W2V121),
				.b6(W2V201),
				.b7(W2V211),
				.b8(W2V221),
				.c(c2100V)
);

ninexnine_unit ninexnine_unit_7430(
				.clk(clk),
				.rstn(rstn),
				.a0(P2002),
				.a1(P2012),
				.a2(P2022),
				.a3(P2102),
				.a4(P2112),
				.a5(P2122),
				.a6(P2202),
				.a7(P2212),
				.a8(P2222),
				.b0(W2V002),
				.b1(W2V012),
				.b2(W2V022),
				.b3(W2V102),
				.b4(W2V112),
				.b5(W2V122),
				.b6(W2V202),
				.b7(W2V212),
				.b8(W2V222),
				.c(c2200V)
);

ninexnine_unit ninexnine_unit_7431(
				.clk(clk),
				.rstn(rstn),
				.a0(P2003),
				.a1(P2013),
				.a2(P2023),
				.a3(P2103),
				.a4(P2113),
				.a5(P2123),
				.a6(P2203),
				.a7(P2213),
				.a8(P2223),
				.b0(W2V003),
				.b1(W2V013),
				.b2(W2V023),
				.b3(W2V103),
				.b4(W2V113),
				.b5(W2V123),
				.b6(W2V203),
				.b7(W2V213),
				.b8(W2V223),
				.c(c2300V)
);

ninexnine_unit ninexnine_unit_7432(
				.clk(clk),
				.rstn(rstn),
				.a0(P2004),
				.a1(P2014),
				.a2(P2024),
				.a3(P2104),
				.a4(P2114),
				.a5(P2124),
				.a6(P2204),
				.a7(P2214),
				.a8(P2224),
				.b0(W2V004),
				.b1(W2V014),
				.b2(W2V024),
				.b3(W2V104),
				.b4(W2V114),
				.b5(W2V124),
				.b6(W2V204),
				.b7(W2V214),
				.b8(W2V224),
				.c(c2400V)
);

ninexnine_unit ninexnine_unit_7433(
				.clk(clk),
				.rstn(rstn),
				.a0(P2005),
				.a1(P2015),
				.a2(P2025),
				.a3(P2105),
				.a4(P2115),
				.a5(P2125),
				.a6(P2205),
				.a7(P2215),
				.a8(P2225),
				.b0(W2V005),
				.b1(W2V015),
				.b2(W2V025),
				.b3(W2V105),
				.b4(W2V115),
				.b5(W2V125),
				.b6(W2V205),
				.b7(W2V215),
				.b8(W2V225),
				.c(c2500V)
);

ninexnine_unit ninexnine_unit_7434(
				.clk(clk),
				.rstn(rstn),
				.a0(P2006),
				.a1(P2016),
				.a2(P2026),
				.a3(P2106),
				.a4(P2116),
				.a5(P2126),
				.a6(P2206),
				.a7(P2216),
				.a8(P2226),
				.b0(W2V006),
				.b1(W2V016),
				.b2(W2V026),
				.b3(W2V106),
				.b4(W2V116),
				.b5(W2V126),
				.b6(W2V206),
				.b7(W2V216),
				.b8(W2V226),
				.c(c2600V)
);

ninexnine_unit ninexnine_unit_7435(
				.clk(clk),
				.rstn(rstn),
				.a0(P2007),
				.a1(P2017),
				.a2(P2027),
				.a3(P2107),
				.a4(P2117),
				.a5(P2127),
				.a6(P2207),
				.a7(P2217),
				.a8(P2227),
				.b0(W2V007),
				.b1(W2V017),
				.b2(W2V027),
				.b3(W2V107),
				.b4(W2V117),
				.b5(W2V127),
				.b6(W2V207),
				.b7(W2V217),
				.b8(W2V227),
				.c(c2700V)
);

ninexnine_unit ninexnine_unit_7436(
				.clk(clk),
				.rstn(rstn),
				.a0(P2008),
				.a1(P2018),
				.a2(P2028),
				.a3(P2108),
				.a4(P2118),
				.a5(P2128),
				.a6(P2208),
				.a7(P2218),
				.a8(P2228),
				.b0(W2V008),
				.b1(W2V018),
				.b2(W2V028),
				.b3(W2V108),
				.b4(W2V118),
				.b5(W2V128),
				.b6(W2V208),
				.b7(W2V218),
				.b8(W2V228),
				.c(c2800V)
);

ninexnine_unit ninexnine_unit_7437(
				.clk(clk),
				.rstn(rstn),
				.a0(P2009),
				.a1(P2019),
				.a2(P2029),
				.a3(P2109),
				.a4(P2119),
				.a5(P2129),
				.a6(P2209),
				.a7(P2219),
				.a8(P2229),
				.b0(W2V009),
				.b1(W2V019),
				.b2(W2V029),
				.b3(W2V109),
				.b4(W2V119),
				.b5(W2V129),
				.b6(W2V209),
				.b7(W2V219),
				.b8(W2V229),
				.c(c2900V)
);

ninexnine_unit ninexnine_unit_7438(
				.clk(clk),
				.rstn(rstn),
				.a0(P200A),
				.a1(P201A),
				.a2(P202A),
				.a3(P210A),
				.a4(P211A),
				.a5(P212A),
				.a6(P220A),
				.a7(P221A),
				.a8(P222A),
				.b0(W2V00A),
				.b1(W2V01A),
				.b2(W2V02A),
				.b3(W2V10A),
				.b4(W2V11A),
				.b5(W2V12A),
				.b6(W2V20A),
				.b7(W2V21A),
				.b8(W2V22A),
				.c(c2A00V)
);

ninexnine_unit ninexnine_unit_7439(
				.clk(clk),
				.rstn(rstn),
				.a0(P200B),
				.a1(P201B),
				.a2(P202B),
				.a3(P210B),
				.a4(P211B),
				.a5(P212B),
				.a6(P220B),
				.a7(P221B),
				.a8(P222B),
				.b0(W2V00B),
				.b1(W2V01B),
				.b2(W2V02B),
				.b3(W2V10B),
				.b4(W2V11B),
				.b5(W2V12B),
				.b6(W2V20B),
				.b7(W2V21B),
				.b8(W2V22B),
				.c(c2B00V)
);

ninexnine_unit ninexnine_unit_7440(
				.clk(clk),
				.rstn(rstn),
				.a0(P200C),
				.a1(P201C),
				.a2(P202C),
				.a3(P210C),
				.a4(P211C),
				.a5(P212C),
				.a6(P220C),
				.a7(P221C),
				.a8(P222C),
				.b0(W2V00C),
				.b1(W2V01C),
				.b2(W2V02C),
				.b3(W2V10C),
				.b4(W2V11C),
				.b5(W2V12C),
				.b6(W2V20C),
				.b7(W2V21C),
				.b8(W2V22C),
				.c(c2C00V)
);

ninexnine_unit ninexnine_unit_7441(
				.clk(clk),
				.rstn(rstn),
				.a0(P200D),
				.a1(P201D),
				.a2(P202D),
				.a3(P210D),
				.a4(P211D),
				.a5(P212D),
				.a6(P220D),
				.a7(P221D),
				.a8(P222D),
				.b0(W2V00D),
				.b1(W2V01D),
				.b2(W2V02D),
				.b3(W2V10D),
				.b4(W2V11D),
				.b5(W2V12D),
				.b6(W2V20D),
				.b7(W2V21D),
				.b8(W2V22D),
				.c(c2D00V)
);

ninexnine_unit ninexnine_unit_7442(
				.clk(clk),
				.rstn(rstn),
				.a0(P200E),
				.a1(P201E),
				.a2(P202E),
				.a3(P210E),
				.a4(P211E),
				.a5(P212E),
				.a6(P220E),
				.a7(P221E),
				.a8(P222E),
				.b0(W2V00E),
				.b1(W2V01E),
				.b2(W2V02E),
				.b3(W2V10E),
				.b4(W2V11E),
				.b5(W2V12E),
				.b6(W2V20E),
				.b7(W2V21E),
				.b8(W2V22E),
				.c(c2E00V)
);

ninexnine_unit ninexnine_unit_7443(
				.clk(clk),
				.rstn(rstn),
				.a0(P200F),
				.a1(P201F),
				.a2(P202F),
				.a3(P210F),
				.a4(P211F),
				.a5(P212F),
				.a6(P220F),
				.a7(P221F),
				.a8(P222F),
				.b0(W2V00F),
				.b1(W2V01F),
				.b2(W2V02F),
				.b3(W2V10F),
				.b4(W2V11F),
				.b5(W2V12F),
				.b6(W2V20F),
				.b7(W2V21F),
				.b8(W2V22F),
				.c(c2F00V)
);

assign C200V=c2000V+c2100V+c2200V+c2300V+c2400V+c2500V+c2600V+c2700V+c2800V+c2900V+c2A00V+c2B00V+c2C00V+c2D00V+c2E00V+c2F00V;
assign A200V=(C200V>=0)?1:0;

assign P300V=A200V;

ninexnine_unit ninexnine_unit_7444(
				.clk(clk),
				.rstn(rstn),
				.a0(P2010),
				.a1(P2020),
				.a2(P2030),
				.a3(P2110),
				.a4(P2120),
				.a5(P2130),
				.a6(P2210),
				.a7(P2220),
				.a8(P2230),
				.b0(W2V000),
				.b1(W2V010),
				.b2(W2V020),
				.b3(W2V100),
				.b4(W2V110),
				.b5(W2V120),
				.b6(W2V200),
				.b7(W2V210),
				.b8(W2V220),
				.c(c2001V)
);

ninexnine_unit ninexnine_unit_7445(
				.clk(clk),
				.rstn(rstn),
				.a0(P2011),
				.a1(P2021),
				.a2(P2031),
				.a3(P2111),
				.a4(P2121),
				.a5(P2131),
				.a6(P2211),
				.a7(P2221),
				.a8(P2231),
				.b0(W2V001),
				.b1(W2V011),
				.b2(W2V021),
				.b3(W2V101),
				.b4(W2V111),
				.b5(W2V121),
				.b6(W2V201),
				.b7(W2V211),
				.b8(W2V221),
				.c(c2101V)
);

ninexnine_unit ninexnine_unit_7446(
				.clk(clk),
				.rstn(rstn),
				.a0(P2012),
				.a1(P2022),
				.a2(P2032),
				.a3(P2112),
				.a4(P2122),
				.a5(P2132),
				.a6(P2212),
				.a7(P2222),
				.a8(P2232),
				.b0(W2V002),
				.b1(W2V012),
				.b2(W2V022),
				.b3(W2V102),
				.b4(W2V112),
				.b5(W2V122),
				.b6(W2V202),
				.b7(W2V212),
				.b8(W2V222),
				.c(c2201V)
);

ninexnine_unit ninexnine_unit_7447(
				.clk(clk),
				.rstn(rstn),
				.a0(P2013),
				.a1(P2023),
				.a2(P2033),
				.a3(P2113),
				.a4(P2123),
				.a5(P2133),
				.a6(P2213),
				.a7(P2223),
				.a8(P2233),
				.b0(W2V003),
				.b1(W2V013),
				.b2(W2V023),
				.b3(W2V103),
				.b4(W2V113),
				.b5(W2V123),
				.b6(W2V203),
				.b7(W2V213),
				.b8(W2V223),
				.c(c2301V)
);

ninexnine_unit ninexnine_unit_7448(
				.clk(clk),
				.rstn(rstn),
				.a0(P2014),
				.a1(P2024),
				.a2(P2034),
				.a3(P2114),
				.a4(P2124),
				.a5(P2134),
				.a6(P2214),
				.a7(P2224),
				.a8(P2234),
				.b0(W2V004),
				.b1(W2V014),
				.b2(W2V024),
				.b3(W2V104),
				.b4(W2V114),
				.b5(W2V124),
				.b6(W2V204),
				.b7(W2V214),
				.b8(W2V224),
				.c(c2401V)
);

ninexnine_unit ninexnine_unit_7449(
				.clk(clk),
				.rstn(rstn),
				.a0(P2015),
				.a1(P2025),
				.a2(P2035),
				.a3(P2115),
				.a4(P2125),
				.a5(P2135),
				.a6(P2215),
				.a7(P2225),
				.a8(P2235),
				.b0(W2V005),
				.b1(W2V015),
				.b2(W2V025),
				.b3(W2V105),
				.b4(W2V115),
				.b5(W2V125),
				.b6(W2V205),
				.b7(W2V215),
				.b8(W2V225),
				.c(c2501V)
);

ninexnine_unit ninexnine_unit_7450(
				.clk(clk),
				.rstn(rstn),
				.a0(P2016),
				.a1(P2026),
				.a2(P2036),
				.a3(P2116),
				.a4(P2126),
				.a5(P2136),
				.a6(P2216),
				.a7(P2226),
				.a8(P2236),
				.b0(W2V006),
				.b1(W2V016),
				.b2(W2V026),
				.b3(W2V106),
				.b4(W2V116),
				.b5(W2V126),
				.b6(W2V206),
				.b7(W2V216),
				.b8(W2V226),
				.c(c2601V)
);

ninexnine_unit ninexnine_unit_7451(
				.clk(clk),
				.rstn(rstn),
				.a0(P2017),
				.a1(P2027),
				.a2(P2037),
				.a3(P2117),
				.a4(P2127),
				.a5(P2137),
				.a6(P2217),
				.a7(P2227),
				.a8(P2237),
				.b0(W2V007),
				.b1(W2V017),
				.b2(W2V027),
				.b3(W2V107),
				.b4(W2V117),
				.b5(W2V127),
				.b6(W2V207),
				.b7(W2V217),
				.b8(W2V227),
				.c(c2701V)
);

ninexnine_unit ninexnine_unit_7452(
				.clk(clk),
				.rstn(rstn),
				.a0(P2018),
				.a1(P2028),
				.a2(P2038),
				.a3(P2118),
				.a4(P2128),
				.a5(P2138),
				.a6(P2218),
				.a7(P2228),
				.a8(P2238),
				.b0(W2V008),
				.b1(W2V018),
				.b2(W2V028),
				.b3(W2V108),
				.b4(W2V118),
				.b5(W2V128),
				.b6(W2V208),
				.b7(W2V218),
				.b8(W2V228),
				.c(c2801V)
);

ninexnine_unit ninexnine_unit_7453(
				.clk(clk),
				.rstn(rstn),
				.a0(P2019),
				.a1(P2029),
				.a2(P2039),
				.a3(P2119),
				.a4(P2129),
				.a5(P2139),
				.a6(P2219),
				.a7(P2229),
				.a8(P2239),
				.b0(W2V009),
				.b1(W2V019),
				.b2(W2V029),
				.b3(W2V109),
				.b4(W2V119),
				.b5(W2V129),
				.b6(W2V209),
				.b7(W2V219),
				.b8(W2V229),
				.c(c2901V)
);

ninexnine_unit ninexnine_unit_7454(
				.clk(clk),
				.rstn(rstn),
				.a0(P201A),
				.a1(P202A),
				.a2(P203A),
				.a3(P211A),
				.a4(P212A),
				.a5(P213A),
				.a6(P221A),
				.a7(P222A),
				.a8(P223A),
				.b0(W2V00A),
				.b1(W2V01A),
				.b2(W2V02A),
				.b3(W2V10A),
				.b4(W2V11A),
				.b5(W2V12A),
				.b6(W2V20A),
				.b7(W2V21A),
				.b8(W2V22A),
				.c(c2A01V)
);

ninexnine_unit ninexnine_unit_7455(
				.clk(clk),
				.rstn(rstn),
				.a0(P201B),
				.a1(P202B),
				.a2(P203B),
				.a3(P211B),
				.a4(P212B),
				.a5(P213B),
				.a6(P221B),
				.a7(P222B),
				.a8(P223B),
				.b0(W2V00B),
				.b1(W2V01B),
				.b2(W2V02B),
				.b3(W2V10B),
				.b4(W2V11B),
				.b5(W2V12B),
				.b6(W2V20B),
				.b7(W2V21B),
				.b8(W2V22B),
				.c(c2B01V)
);

ninexnine_unit ninexnine_unit_7456(
				.clk(clk),
				.rstn(rstn),
				.a0(P201C),
				.a1(P202C),
				.a2(P203C),
				.a3(P211C),
				.a4(P212C),
				.a5(P213C),
				.a6(P221C),
				.a7(P222C),
				.a8(P223C),
				.b0(W2V00C),
				.b1(W2V01C),
				.b2(W2V02C),
				.b3(W2V10C),
				.b4(W2V11C),
				.b5(W2V12C),
				.b6(W2V20C),
				.b7(W2V21C),
				.b8(W2V22C),
				.c(c2C01V)
);

ninexnine_unit ninexnine_unit_7457(
				.clk(clk),
				.rstn(rstn),
				.a0(P201D),
				.a1(P202D),
				.a2(P203D),
				.a3(P211D),
				.a4(P212D),
				.a5(P213D),
				.a6(P221D),
				.a7(P222D),
				.a8(P223D),
				.b0(W2V00D),
				.b1(W2V01D),
				.b2(W2V02D),
				.b3(W2V10D),
				.b4(W2V11D),
				.b5(W2V12D),
				.b6(W2V20D),
				.b7(W2V21D),
				.b8(W2V22D),
				.c(c2D01V)
);

ninexnine_unit ninexnine_unit_7458(
				.clk(clk),
				.rstn(rstn),
				.a0(P201E),
				.a1(P202E),
				.a2(P203E),
				.a3(P211E),
				.a4(P212E),
				.a5(P213E),
				.a6(P221E),
				.a7(P222E),
				.a8(P223E),
				.b0(W2V00E),
				.b1(W2V01E),
				.b2(W2V02E),
				.b3(W2V10E),
				.b4(W2V11E),
				.b5(W2V12E),
				.b6(W2V20E),
				.b7(W2V21E),
				.b8(W2V22E),
				.c(c2E01V)
);

ninexnine_unit ninexnine_unit_7459(
				.clk(clk),
				.rstn(rstn),
				.a0(P201F),
				.a1(P202F),
				.a2(P203F),
				.a3(P211F),
				.a4(P212F),
				.a5(P213F),
				.a6(P221F),
				.a7(P222F),
				.a8(P223F),
				.b0(W2V00F),
				.b1(W2V01F),
				.b2(W2V02F),
				.b3(W2V10F),
				.b4(W2V11F),
				.b5(W2V12F),
				.b6(W2V20F),
				.b7(W2V21F),
				.b8(W2V22F),
				.c(c2F01V)
);

assign C201V=c2001V+c2101V+c2201V+c2301V+c2401V+c2501V+c2601V+c2701V+c2801V+c2901V+c2A01V+c2B01V+c2C01V+c2D01V+c2E01V+c2F01V;
assign A201V=(C201V>=0)?1:0;

assign P301V=A201V;

ninexnine_unit ninexnine_unit_7460(
				.clk(clk),
				.rstn(rstn),
				.a0(P2020),
				.a1(P2030),
				.a2(P2040),
				.a3(P2120),
				.a4(P2130),
				.a5(P2140),
				.a6(P2220),
				.a7(P2230),
				.a8(P2240),
				.b0(W2V000),
				.b1(W2V010),
				.b2(W2V020),
				.b3(W2V100),
				.b4(W2V110),
				.b5(W2V120),
				.b6(W2V200),
				.b7(W2V210),
				.b8(W2V220),
				.c(c2002V)
);

ninexnine_unit ninexnine_unit_7461(
				.clk(clk),
				.rstn(rstn),
				.a0(P2021),
				.a1(P2031),
				.a2(P2041),
				.a3(P2121),
				.a4(P2131),
				.a5(P2141),
				.a6(P2221),
				.a7(P2231),
				.a8(P2241),
				.b0(W2V001),
				.b1(W2V011),
				.b2(W2V021),
				.b3(W2V101),
				.b4(W2V111),
				.b5(W2V121),
				.b6(W2V201),
				.b7(W2V211),
				.b8(W2V221),
				.c(c2102V)
);

ninexnine_unit ninexnine_unit_7462(
				.clk(clk),
				.rstn(rstn),
				.a0(P2022),
				.a1(P2032),
				.a2(P2042),
				.a3(P2122),
				.a4(P2132),
				.a5(P2142),
				.a6(P2222),
				.a7(P2232),
				.a8(P2242),
				.b0(W2V002),
				.b1(W2V012),
				.b2(W2V022),
				.b3(W2V102),
				.b4(W2V112),
				.b5(W2V122),
				.b6(W2V202),
				.b7(W2V212),
				.b8(W2V222),
				.c(c2202V)
);

ninexnine_unit ninexnine_unit_7463(
				.clk(clk),
				.rstn(rstn),
				.a0(P2023),
				.a1(P2033),
				.a2(P2043),
				.a3(P2123),
				.a4(P2133),
				.a5(P2143),
				.a6(P2223),
				.a7(P2233),
				.a8(P2243),
				.b0(W2V003),
				.b1(W2V013),
				.b2(W2V023),
				.b3(W2V103),
				.b4(W2V113),
				.b5(W2V123),
				.b6(W2V203),
				.b7(W2V213),
				.b8(W2V223),
				.c(c2302V)
);

ninexnine_unit ninexnine_unit_7464(
				.clk(clk),
				.rstn(rstn),
				.a0(P2024),
				.a1(P2034),
				.a2(P2044),
				.a3(P2124),
				.a4(P2134),
				.a5(P2144),
				.a6(P2224),
				.a7(P2234),
				.a8(P2244),
				.b0(W2V004),
				.b1(W2V014),
				.b2(W2V024),
				.b3(W2V104),
				.b4(W2V114),
				.b5(W2V124),
				.b6(W2V204),
				.b7(W2V214),
				.b8(W2V224),
				.c(c2402V)
);

ninexnine_unit ninexnine_unit_7465(
				.clk(clk),
				.rstn(rstn),
				.a0(P2025),
				.a1(P2035),
				.a2(P2045),
				.a3(P2125),
				.a4(P2135),
				.a5(P2145),
				.a6(P2225),
				.a7(P2235),
				.a8(P2245),
				.b0(W2V005),
				.b1(W2V015),
				.b2(W2V025),
				.b3(W2V105),
				.b4(W2V115),
				.b5(W2V125),
				.b6(W2V205),
				.b7(W2V215),
				.b8(W2V225),
				.c(c2502V)
);

ninexnine_unit ninexnine_unit_7466(
				.clk(clk),
				.rstn(rstn),
				.a0(P2026),
				.a1(P2036),
				.a2(P2046),
				.a3(P2126),
				.a4(P2136),
				.a5(P2146),
				.a6(P2226),
				.a7(P2236),
				.a8(P2246),
				.b0(W2V006),
				.b1(W2V016),
				.b2(W2V026),
				.b3(W2V106),
				.b4(W2V116),
				.b5(W2V126),
				.b6(W2V206),
				.b7(W2V216),
				.b8(W2V226),
				.c(c2602V)
);

ninexnine_unit ninexnine_unit_7467(
				.clk(clk),
				.rstn(rstn),
				.a0(P2027),
				.a1(P2037),
				.a2(P2047),
				.a3(P2127),
				.a4(P2137),
				.a5(P2147),
				.a6(P2227),
				.a7(P2237),
				.a8(P2247),
				.b0(W2V007),
				.b1(W2V017),
				.b2(W2V027),
				.b3(W2V107),
				.b4(W2V117),
				.b5(W2V127),
				.b6(W2V207),
				.b7(W2V217),
				.b8(W2V227),
				.c(c2702V)
);

ninexnine_unit ninexnine_unit_7468(
				.clk(clk),
				.rstn(rstn),
				.a0(P2028),
				.a1(P2038),
				.a2(P2048),
				.a3(P2128),
				.a4(P2138),
				.a5(P2148),
				.a6(P2228),
				.a7(P2238),
				.a8(P2248),
				.b0(W2V008),
				.b1(W2V018),
				.b2(W2V028),
				.b3(W2V108),
				.b4(W2V118),
				.b5(W2V128),
				.b6(W2V208),
				.b7(W2V218),
				.b8(W2V228),
				.c(c2802V)
);

ninexnine_unit ninexnine_unit_7469(
				.clk(clk),
				.rstn(rstn),
				.a0(P2029),
				.a1(P2039),
				.a2(P2049),
				.a3(P2129),
				.a4(P2139),
				.a5(P2149),
				.a6(P2229),
				.a7(P2239),
				.a8(P2249),
				.b0(W2V009),
				.b1(W2V019),
				.b2(W2V029),
				.b3(W2V109),
				.b4(W2V119),
				.b5(W2V129),
				.b6(W2V209),
				.b7(W2V219),
				.b8(W2V229),
				.c(c2902V)
);

ninexnine_unit ninexnine_unit_7470(
				.clk(clk),
				.rstn(rstn),
				.a0(P202A),
				.a1(P203A),
				.a2(P204A),
				.a3(P212A),
				.a4(P213A),
				.a5(P214A),
				.a6(P222A),
				.a7(P223A),
				.a8(P224A),
				.b0(W2V00A),
				.b1(W2V01A),
				.b2(W2V02A),
				.b3(W2V10A),
				.b4(W2V11A),
				.b5(W2V12A),
				.b6(W2V20A),
				.b7(W2V21A),
				.b8(W2V22A),
				.c(c2A02V)
);

ninexnine_unit ninexnine_unit_7471(
				.clk(clk),
				.rstn(rstn),
				.a0(P202B),
				.a1(P203B),
				.a2(P204B),
				.a3(P212B),
				.a4(P213B),
				.a5(P214B),
				.a6(P222B),
				.a7(P223B),
				.a8(P224B),
				.b0(W2V00B),
				.b1(W2V01B),
				.b2(W2V02B),
				.b3(W2V10B),
				.b4(W2V11B),
				.b5(W2V12B),
				.b6(W2V20B),
				.b7(W2V21B),
				.b8(W2V22B),
				.c(c2B02V)
);

ninexnine_unit ninexnine_unit_7472(
				.clk(clk),
				.rstn(rstn),
				.a0(P202C),
				.a1(P203C),
				.a2(P204C),
				.a3(P212C),
				.a4(P213C),
				.a5(P214C),
				.a6(P222C),
				.a7(P223C),
				.a8(P224C),
				.b0(W2V00C),
				.b1(W2V01C),
				.b2(W2V02C),
				.b3(W2V10C),
				.b4(W2V11C),
				.b5(W2V12C),
				.b6(W2V20C),
				.b7(W2V21C),
				.b8(W2V22C),
				.c(c2C02V)
);

ninexnine_unit ninexnine_unit_7473(
				.clk(clk),
				.rstn(rstn),
				.a0(P202D),
				.a1(P203D),
				.a2(P204D),
				.a3(P212D),
				.a4(P213D),
				.a5(P214D),
				.a6(P222D),
				.a7(P223D),
				.a8(P224D),
				.b0(W2V00D),
				.b1(W2V01D),
				.b2(W2V02D),
				.b3(W2V10D),
				.b4(W2V11D),
				.b5(W2V12D),
				.b6(W2V20D),
				.b7(W2V21D),
				.b8(W2V22D),
				.c(c2D02V)
);

ninexnine_unit ninexnine_unit_7474(
				.clk(clk),
				.rstn(rstn),
				.a0(P202E),
				.a1(P203E),
				.a2(P204E),
				.a3(P212E),
				.a4(P213E),
				.a5(P214E),
				.a6(P222E),
				.a7(P223E),
				.a8(P224E),
				.b0(W2V00E),
				.b1(W2V01E),
				.b2(W2V02E),
				.b3(W2V10E),
				.b4(W2V11E),
				.b5(W2V12E),
				.b6(W2V20E),
				.b7(W2V21E),
				.b8(W2V22E),
				.c(c2E02V)
);

ninexnine_unit ninexnine_unit_7475(
				.clk(clk),
				.rstn(rstn),
				.a0(P202F),
				.a1(P203F),
				.a2(P204F),
				.a3(P212F),
				.a4(P213F),
				.a5(P214F),
				.a6(P222F),
				.a7(P223F),
				.a8(P224F),
				.b0(W2V00F),
				.b1(W2V01F),
				.b2(W2V02F),
				.b3(W2V10F),
				.b4(W2V11F),
				.b5(W2V12F),
				.b6(W2V20F),
				.b7(W2V21F),
				.b8(W2V22F),
				.c(c2F02V)
);

assign C202V=c2002V+c2102V+c2202V+c2302V+c2402V+c2502V+c2602V+c2702V+c2802V+c2902V+c2A02V+c2B02V+c2C02V+c2D02V+c2E02V+c2F02V;
assign A202V=(C202V>=0)?1:0;

assign P302V=A202V;

ninexnine_unit ninexnine_unit_7476(
				.clk(clk),
				.rstn(rstn),
				.a0(P2100),
				.a1(P2110),
				.a2(P2120),
				.a3(P2200),
				.a4(P2210),
				.a5(P2220),
				.a6(P2300),
				.a7(P2310),
				.a8(P2320),
				.b0(W2V000),
				.b1(W2V010),
				.b2(W2V020),
				.b3(W2V100),
				.b4(W2V110),
				.b5(W2V120),
				.b6(W2V200),
				.b7(W2V210),
				.b8(W2V220),
				.c(c2010V)
);

ninexnine_unit ninexnine_unit_7477(
				.clk(clk),
				.rstn(rstn),
				.a0(P2101),
				.a1(P2111),
				.a2(P2121),
				.a3(P2201),
				.a4(P2211),
				.a5(P2221),
				.a6(P2301),
				.a7(P2311),
				.a8(P2321),
				.b0(W2V001),
				.b1(W2V011),
				.b2(W2V021),
				.b3(W2V101),
				.b4(W2V111),
				.b5(W2V121),
				.b6(W2V201),
				.b7(W2V211),
				.b8(W2V221),
				.c(c2110V)
);

ninexnine_unit ninexnine_unit_7478(
				.clk(clk),
				.rstn(rstn),
				.a0(P2102),
				.a1(P2112),
				.a2(P2122),
				.a3(P2202),
				.a4(P2212),
				.a5(P2222),
				.a6(P2302),
				.a7(P2312),
				.a8(P2322),
				.b0(W2V002),
				.b1(W2V012),
				.b2(W2V022),
				.b3(W2V102),
				.b4(W2V112),
				.b5(W2V122),
				.b6(W2V202),
				.b7(W2V212),
				.b8(W2V222),
				.c(c2210V)
);

ninexnine_unit ninexnine_unit_7479(
				.clk(clk),
				.rstn(rstn),
				.a0(P2103),
				.a1(P2113),
				.a2(P2123),
				.a3(P2203),
				.a4(P2213),
				.a5(P2223),
				.a6(P2303),
				.a7(P2313),
				.a8(P2323),
				.b0(W2V003),
				.b1(W2V013),
				.b2(W2V023),
				.b3(W2V103),
				.b4(W2V113),
				.b5(W2V123),
				.b6(W2V203),
				.b7(W2V213),
				.b8(W2V223),
				.c(c2310V)
);

ninexnine_unit ninexnine_unit_7480(
				.clk(clk),
				.rstn(rstn),
				.a0(P2104),
				.a1(P2114),
				.a2(P2124),
				.a3(P2204),
				.a4(P2214),
				.a5(P2224),
				.a6(P2304),
				.a7(P2314),
				.a8(P2324),
				.b0(W2V004),
				.b1(W2V014),
				.b2(W2V024),
				.b3(W2V104),
				.b4(W2V114),
				.b5(W2V124),
				.b6(W2V204),
				.b7(W2V214),
				.b8(W2V224),
				.c(c2410V)
);

ninexnine_unit ninexnine_unit_7481(
				.clk(clk),
				.rstn(rstn),
				.a0(P2105),
				.a1(P2115),
				.a2(P2125),
				.a3(P2205),
				.a4(P2215),
				.a5(P2225),
				.a6(P2305),
				.a7(P2315),
				.a8(P2325),
				.b0(W2V005),
				.b1(W2V015),
				.b2(W2V025),
				.b3(W2V105),
				.b4(W2V115),
				.b5(W2V125),
				.b6(W2V205),
				.b7(W2V215),
				.b8(W2V225),
				.c(c2510V)
);

ninexnine_unit ninexnine_unit_7482(
				.clk(clk),
				.rstn(rstn),
				.a0(P2106),
				.a1(P2116),
				.a2(P2126),
				.a3(P2206),
				.a4(P2216),
				.a5(P2226),
				.a6(P2306),
				.a7(P2316),
				.a8(P2326),
				.b0(W2V006),
				.b1(W2V016),
				.b2(W2V026),
				.b3(W2V106),
				.b4(W2V116),
				.b5(W2V126),
				.b6(W2V206),
				.b7(W2V216),
				.b8(W2V226),
				.c(c2610V)
);

ninexnine_unit ninexnine_unit_7483(
				.clk(clk),
				.rstn(rstn),
				.a0(P2107),
				.a1(P2117),
				.a2(P2127),
				.a3(P2207),
				.a4(P2217),
				.a5(P2227),
				.a6(P2307),
				.a7(P2317),
				.a8(P2327),
				.b0(W2V007),
				.b1(W2V017),
				.b2(W2V027),
				.b3(W2V107),
				.b4(W2V117),
				.b5(W2V127),
				.b6(W2V207),
				.b7(W2V217),
				.b8(W2V227),
				.c(c2710V)
);

ninexnine_unit ninexnine_unit_7484(
				.clk(clk),
				.rstn(rstn),
				.a0(P2108),
				.a1(P2118),
				.a2(P2128),
				.a3(P2208),
				.a4(P2218),
				.a5(P2228),
				.a6(P2308),
				.a7(P2318),
				.a8(P2328),
				.b0(W2V008),
				.b1(W2V018),
				.b2(W2V028),
				.b3(W2V108),
				.b4(W2V118),
				.b5(W2V128),
				.b6(W2V208),
				.b7(W2V218),
				.b8(W2V228),
				.c(c2810V)
);

ninexnine_unit ninexnine_unit_7485(
				.clk(clk),
				.rstn(rstn),
				.a0(P2109),
				.a1(P2119),
				.a2(P2129),
				.a3(P2209),
				.a4(P2219),
				.a5(P2229),
				.a6(P2309),
				.a7(P2319),
				.a8(P2329),
				.b0(W2V009),
				.b1(W2V019),
				.b2(W2V029),
				.b3(W2V109),
				.b4(W2V119),
				.b5(W2V129),
				.b6(W2V209),
				.b7(W2V219),
				.b8(W2V229),
				.c(c2910V)
);

ninexnine_unit ninexnine_unit_7486(
				.clk(clk),
				.rstn(rstn),
				.a0(P210A),
				.a1(P211A),
				.a2(P212A),
				.a3(P220A),
				.a4(P221A),
				.a5(P222A),
				.a6(P230A),
				.a7(P231A),
				.a8(P232A),
				.b0(W2V00A),
				.b1(W2V01A),
				.b2(W2V02A),
				.b3(W2V10A),
				.b4(W2V11A),
				.b5(W2V12A),
				.b6(W2V20A),
				.b7(W2V21A),
				.b8(W2V22A),
				.c(c2A10V)
);

ninexnine_unit ninexnine_unit_7487(
				.clk(clk),
				.rstn(rstn),
				.a0(P210B),
				.a1(P211B),
				.a2(P212B),
				.a3(P220B),
				.a4(P221B),
				.a5(P222B),
				.a6(P230B),
				.a7(P231B),
				.a8(P232B),
				.b0(W2V00B),
				.b1(W2V01B),
				.b2(W2V02B),
				.b3(W2V10B),
				.b4(W2V11B),
				.b5(W2V12B),
				.b6(W2V20B),
				.b7(W2V21B),
				.b8(W2V22B),
				.c(c2B10V)
);

ninexnine_unit ninexnine_unit_7488(
				.clk(clk),
				.rstn(rstn),
				.a0(P210C),
				.a1(P211C),
				.a2(P212C),
				.a3(P220C),
				.a4(P221C),
				.a5(P222C),
				.a6(P230C),
				.a7(P231C),
				.a8(P232C),
				.b0(W2V00C),
				.b1(W2V01C),
				.b2(W2V02C),
				.b3(W2V10C),
				.b4(W2V11C),
				.b5(W2V12C),
				.b6(W2V20C),
				.b7(W2V21C),
				.b8(W2V22C),
				.c(c2C10V)
);

ninexnine_unit ninexnine_unit_7489(
				.clk(clk),
				.rstn(rstn),
				.a0(P210D),
				.a1(P211D),
				.a2(P212D),
				.a3(P220D),
				.a4(P221D),
				.a5(P222D),
				.a6(P230D),
				.a7(P231D),
				.a8(P232D),
				.b0(W2V00D),
				.b1(W2V01D),
				.b2(W2V02D),
				.b3(W2V10D),
				.b4(W2V11D),
				.b5(W2V12D),
				.b6(W2V20D),
				.b7(W2V21D),
				.b8(W2V22D),
				.c(c2D10V)
);

ninexnine_unit ninexnine_unit_7490(
				.clk(clk),
				.rstn(rstn),
				.a0(P210E),
				.a1(P211E),
				.a2(P212E),
				.a3(P220E),
				.a4(P221E),
				.a5(P222E),
				.a6(P230E),
				.a7(P231E),
				.a8(P232E),
				.b0(W2V00E),
				.b1(W2V01E),
				.b2(W2V02E),
				.b3(W2V10E),
				.b4(W2V11E),
				.b5(W2V12E),
				.b6(W2V20E),
				.b7(W2V21E),
				.b8(W2V22E),
				.c(c2E10V)
);

ninexnine_unit ninexnine_unit_7491(
				.clk(clk),
				.rstn(rstn),
				.a0(P210F),
				.a1(P211F),
				.a2(P212F),
				.a3(P220F),
				.a4(P221F),
				.a5(P222F),
				.a6(P230F),
				.a7(P231F),
				.a8(P232F),
				.b0(W2V00F),
				.b1(W2V01F),
				.b2(W2V02F),
				.b3(W2V10F),
				.b4(W2V11F),
				.b5(W2V12F),
				.b6(W2V20F),
				.b7(W2V21F),
				.b8(W2V22F),
				.c(c2F10V)
);

assign C210V=c2010V+c2110V+c2210V+c2310V+c2410V+c2510V+c2610V+c2710V+c2810V+c2910V+c2A10V+c2B10V+c2C10V+c2D10V+c2E10V+c2F10V;
assign A210V=(C210V>=0)?1:0;

assign P310V=A210V;

ninexnine_unit ninexnine_unit_7492(
				.clk(clk),
				.rstn(rstn),
				.a0(P2110),
				.a1(P2120),
				.a2(P2130),
				.a3(P2210),
				.a4(P2220),
				.a5(P2230),
				.a6(P2310),
				.a7(P2320),
				.a8(P2330),
				.b0(W2V000),
				.b1(W2V010),
				.b2(W2V020),
				.b3(W2V100),
				.b4(W2V110),
				.b5(W2V120),
				.b6(W2V200),
				.b7(W2V210),
				.b8(W2V220),
				.c(c2011V)
);

ninexnine_unit ninexnine_unit_7493(
				.clk(clk),
				.rstn(rstn),
				.a0(P2111),
				.a1(P2121),
				.a2(P2131),
				.a3(P2211),
				.a4(P2221),
				.a5(P2231),
				.a6(P2311),
				.a7(P2321),
				.a8(P2331),
				.b0(W2V001),
				.b1(W2V011),
				.b2(W2V021),
				.b3(W2V101),
				.b4(W2V111),
				.b5(W2V121),
				.b6(W2V201),
				.b7(W2V211),
				.b8(W2V221),
				.c(c2111V)
);

ninexnine_unit ninexnine_unit_7494(
				.clk(clk),
				.rstn(rstn),
				.a0(P2112),
				.a1(P2122),
				.a2(P2132),
				.a3(P2212),
				.a4(P2222),
				.a5(P2232),
				.a6(P2312),
				.a7(P2322),
				.a8(P2332),
				.b0(W2V002),
				.b1(W2V012),
				.b2(W2V022),
				.b3(W2V102),
				.b4(W2V112),
				.b5(W2V122),
				.b6(W2V202),
				.b7(W2V212),
				.b8(W2V222),
				.c(c2211V)
);

ninexnine_unit ninexnine_unit_7495(
				.clk(clk),
				.rstn(rstn),
				.a0(P2113),
				.a1(P2123),
				.a2(P2133),
				.a3(P2213),
				.a4(P2223),
				.a5(P2233),
				.a6(P2313),
				.a7(P2323),
				.a8(P2333),
				.b0(W2V003),
				.b1(W2V013),
				.b2(W2V023),
				.b3(W2V103),
				.b4(W2V113),
				.b5(W2V123),
				.b6(W2V203),
				.b7(W2V213),
				.b8(W2V223),
				.c(c2311V)
);

ninexnine_unit ninexnine_unit_7496(
				.clk(clk),
				.rstn(rstn),
				.a0(P2114),
				.a1(P2124),
				.a2(P2134),
				.a3(P2214),
				.a4(P2224),
				.a5(P2234),
				.a6(P2314),
				.a7(P2324),
				.a8(P2334),
				.b0(W2V004),
				.b1(W2V014),
				.b2(W2V024),
				.b3(W2V104),
				.b4(W2V114),
				.b5(W2V124),
				.b6(W2V204),
				.b7(W2V214),
				.b8(W2V224),
				.c(c2411V)
);

ninexnine_unit ninexnine_unit_7497(
				.clk(clk),
				.rstn(rstn),
				.a0(P2115),
				.a1(P2125),
				.a2(P2135),
				.a3(P2215),
				.a4(P2225),
				.a5(P2235),
				.a6(P2315),
				.a7(P2325),
				.a8(P2335),
				.b0(W2V005),
				.b1(W2V015),
				.b2(W2V025),
				.b3(W2V105),
				.b4(W2V115),
				.b5(W2V125),
				.b6(W2V205),
				.b7(W2V215),
				.b8(W2V225),
				.c(c2511V)
);

ninexnine_unit ninexnine_unit_7498(
				.clk(clk),
				.rstn(rstn),
				.a0(P2116),
				.a1(P2126),
				.a2(P2136),
				.a3(P2216),
				.a4(P2226),
				.a5(P2236),
				.a6(P2316),
				.a7(P2326),
				.a8(P2336),
				.b0(W2V006),
				.b1(W2V016),
				.b2(W2V026),
				.b3(W2V106),
				.b4(W2V116),
				.b5(W2V126),
				.b6(W2V206),
				.b7(W2V216),
				.b8(W2V226),
				.c(c2611V)
);

ninexnine_unit ninexnine_unit_7499(
				.clk(clk),
				.rstn(rstn),
				.a0(P2117),
				.a1(P2127),
				.a2(P2137),
				.a3(P2217),
				.a4(P2227),
				.a5(P2237),
				.a6(P2317),
				.a7(P2327),
				.a8(P2337),
				.b0(W2V007),
				.b1(W2V017),
				.b2(W2V027),
				.b3(W2V107),
				.b4(W2V117),
				.b5(W2V127),
				.b6(W2V207),
				.b7(W2V217),
				.b8(W2V227),
				.c(c2711V)
);

ninexnine_unit ninexnine_unit_7500(
				.clk(clk),
				.rstn(rstn),
				.a0(P2118),
				.a1(P2128),
				.a2(P2138),
				.a3(P2218),
				.a4(P2228),
				.a5(P2238),
				.a6(P2318),
				.a7(P2328),
				.a8(P2338),
				.b0(W2V008),
				.b1(W2V018),
				.b2(W2V028),
				.b3(W2V108),
				.b4(W2V118),
				.b5(W2V128),
				.b6(W2V208),
				.b7(W2V218),
				.b8(W2V228),
				.c(c2811V)
);

ninexnine_unit ninexnine_unit_7501(
				.clk(clk),
				.rstn(rstn),
				.a0(P2119),
				.a1(P2129),
				.a2(P2139),
				.a3(P2219),
				.a4(P2229),
				.a5(P2239),
				.a6(P2319),
				.a7(P2329),
				.a8(P2339),
				.b0(W2V009),
				.b1(W2V019),
				.b2(W2V029),
				.b3(W2V109),
				.b4(W2V119),
				.b5(W2V129),
				.b6(W2V209),
				.b7(W2V219),
				.b8(W2V229),
				.c(c2911V)
);

ninexnine_unit ninexnine_unit_7502(
				.clk(clk),
				.rstn(rstn),
				.a0(P211A),
				.a1(P212A),
				.a2(P213A),
				.a3(P221A),
				.a4(P222A),
				.a5(P223A),
				.a6(P231A),
				.a7(P232A),
				.a8(P233A),
				.b0(W2V00A),
				.b1(W2V01A),
				.b2(W2V02A),
				.b3(W2V10A),
				.b4(W2V11A),
				.b5(W2V12A),
				.b6(W2V20A),
				.b7(W2V21A),
				.b8(W2V22A),
				.c(c2A11V)
);

ninexnine_unit ninexnine_unit_7503(
				.clk(clk),
				.rstn(rstn),
				.a0(P211B),
				.a1(P212B),
				.a2(P213B),
				.a3(P221B),
				.a4(P222B),
				.a5(P223B),
				.a6(P231B),
				.a7(P232B),
				.a8(P233B),
				.b0(W2V00B),
				.b1(W2V01B),
				.b2(W2V02B),
				.b3(W2V10B),
				.b4(W2V11B),
				.b5(W2V12B),
				.b6(W2V20B),
				.b7(W2V21B),
				.b8(W2V22B),
				.c(c2B11V)
);

ninexnine_unit ninexnine_unit_7504(
				.clk(clk),
				.rstn(rstn),
				.a0(P211C),
				.a1(P212C),
				.a2(P213C),
				.a3(P221C),
				.a4(P222C),
				.a5(P223C),
				.a6(P231C),
				.a7(P232C),
				.a8(P233C),
				.b0(W2V00C),
				.b1(W2V01C),
				.b2(W2V02C),
				.b3(W2V10C),
				.b4(W2V11C),
				.b5(W2V12C),
				.b6(W2V20C),
				.b7(W2V21C),
				.b8(W2V22C),
				.c(c2C11V)
);

ninexnine_unit ninexnine_unit_7505(
				.clk(clk),
				.rstn(rstn),
				.a0(P211D),
				.a1(P212D),
				.a2(P213D),
				.a3(P221D),
				.a4(P222D),
				.a5(P223D),
				.a6(P231D),
				.a7(P232D),
				.a8(P233D),
				.b0(W2V00D),
				.b1(W2V01D),
				.b2(W2V02D),
				.b3(W2V10D),
				.b4(W2V11D),
				.b5(W2V12D),
				.b6(W2V20D),
				.b7(W2V21D),
				.b8(W2V22D),
				.c(c2D11V)
);

ninexnine_unit ninexnine_unit_7506(
				.clk(clk),
				.rstn(rstn),
				.a0(P211E),
				.a1(P212E),
				.a2(P213E),
				.a3(P221E),
				.a4(P222E),
				.a5(P223E),
				.a6(P231E),
				.a7(P232E),
				.a8(P233E),
				.b0(W2V00E),
				.b1(W2V01E),
				.b2(W2V02E),
				.b3(W2V10E),
				.b4(W2V11E),
				.b5(W2V12E),
				.b6(W2V20E),
				.b7(W2V21E),
				.b8(W2V22E),
				.c(c2E11V)
);

ninexnine_unit ninexnine_unit_7507(
				.clk(clk),
				.rstn(rstn),
				.a0(P211F),
				.a1(P212F),
				.a2(P213F),
				.a3(P221F),
				.a4(P222F),
				.a5(P223F),
				.a6(P231F),
				.a7(P232F),
				.a8(P233F),
				.b0(W2V00F),
				.b1(W2V01F),
				.b2(W2V02F),
				.b3(W2V10F),
				.b4(W2V11F),
				.b5(W2V12F),
				.b6(W2V20F),
				.b7(W2V21F),
				.b8(W2V22F),
				.c(c2F11V)
);

assign C211V=c2011V+c2111V+c2211V+c2311V+c2411V+c2511V+c2611V+c2711V+c2811V+c2911V+c2A11V+c2B11V+c2C11V+c2D11V+c2E11V+c2F11V;
assign A211V=(C211V>=0)?1:0;

assign P311V=A211V;

ninexnine_unit ninexnine_unit_7508(
				.clk(clk),
				.rstn(rstn),
				.a0(P2120),
				.a1(P2130),
				.a2(P2140),
				.a3(P2220),
				.a4(P2230),
				.a5(P2240),
				.a6(P2320),
				.a7(P2330),
				.a8(P2340),
				.b0(W2V000),
				.b1(W2V010),
				.b2(W2V020),
				.b3(W2V100),
				.b4(W2V110),
				.b5(W2V120),
				.b6(W2V200),
				.b7(W2V210),
				.b8(W2V220),
				.c(c2012V)
);

ninexnine_unit ninexnine_unit_7509(
				.clk(clk),
				.rstn(rstn),
				.a0(P2121),
				.a1(P2131),
				.a2(P2141),
				.a3(P2221),
				.a4(P2231),
				.a5(P2241),
				.a6(P2321),
				.a7(P2331),
				.a8(P2341),
				.b0(W2V001),
				.b1(W2V011),
				.b2(W2V021),
				.b3(W2V101),
				.b4(W2V111),
				.b5(W2V121),
				.b6(W2V201),
				.b7(W2V211),
				.b8(W2V221),
				.c(c2112V)
);

ninexnine_unit ninexnine_unit_7510(
				.clk(clk),
				.rstn(rstn),
				.a0(P2122),
				.a1(P2132),
				.a2(P2142),
				.a3(P2222),
				.a4(P2232),
				.a5(P2242),
				.a6(P2322),
				.a7(P2332),
				.a8(P2342),
				.b0(W2V002),
				.b1(W2V012),
				.b2(W2V022),
				.b3(W2V102),
				.b4(W2V112),
				.b5(W2V122),
				.b6(W2V202),
				.b7(W2V212),
				.b8(W2V222),
				.c(c2212V)
);

ninexnine_unit ninexnine_unit_7511(
				.clk(clk),
				.rstn(rstn),
				.a0(P2123),
				.a1(P2133),
				.a2(P2143),
				.a3(P2223),
				.a4(P2233),
				.a5(P2243),
				.a6(P2323),
				.a7(P2333),
				.a8(P2343),
				.b0(W2V003),
				.b1(W2V013),
				.b2(W2V023),
				.b3(W2V103),
				.b4(W2V113),
				.b5(W2V123),
				.b6(W2V203),
				.b7(W2V213),
				.b8(W2V223),
				.c(c2312V)
);

ninexnine_unit ninexnine_unit_7512(
				.clk(clk),
				.rstn(rstn),
				.a0(P2124),
				.a1(P2134),
				.a2(P2144),
				.a3(P2224),
				.a4(P2234),
				.a5(P2244),
				.a6(P2324),
				.a7(P2334),
				.a8(P2344),
				.b0(W2V004),
				.b1(W2V014),
				.b2(W2V024),
				.b3(W2V104),
				.b4(W2V114),
				.b5(W2V124),
				.b6(W2V204),
				.b7(W2V214),
				.b8(W2V224),
				.c(c2412V)
);

ninexnine_unit ninexnine_unit_7513(
				.clk(clk),
				.rstn(rstn),
				.a0(P2125),
				.a1(P2135),
				.a2(P2145),
				.a3(P2225),
				.a4(P2235),
				.a5(P2245),
				.a6(P2325),
				.a7(P2335),
				.a8(P2345),
				.b0(W2V005),
				.b1(W2V015),
				.b2(W2V025),
				.b3(W2V105),
				.b4(W2V115),
				.b5(W2V125),
				.b6(W2V205),
				.b7(W2V215),
				.b8(W2V225),
				.c(c2512V)
);

ninexnine_unit ninexnine_unit_7514(
				.clk(clk),
				.rstn(rstn),
				.a0(P2126),
				.a1(P2136),
				.a2(P2146),
				.a3(P2226),
				.a4(P2236),
				.a5(P2246),
				.a6(P2326),
				.a7(P2336),
				.a8(P2346),
				.b0(W2V006),
				.b1(W2V016),
				.b2(W2V026),
				.b3(W2V106),
				.b4(W2V116),
				.b5(W2V126),
				.b6(W2V206),
				.b7(W2V216),
				.b8(W2V226),
				.c(c2612V)
);

ninexnine_unit ninexnine_unit_7515(
				.clk(clk),
				.rstn(rstn),
				.a0(P2127),
				.a1(P2137),
				.a2(P2147),
				.a3(P2227),
				.a4(P2237),
				.a5(P2247),
				.a6(P2327),
				.a7(P2337),
				.a8(P2347),
				.b0(W2V007),
				.b1(W2V017),
				.b2(W2V027),
				.b3(W2V107),
				.b4(W2V117),
				.b5(W2V127),
				.b6(W2V207),
				.b7(W2V217),
				.b8(W2V227),
				.c(c2712V)
);

ninexnine_unit ninexnine_unit_7516(
				.clk(clk),
				.rstn(rstn),
				.a0(P2128),
				.a1(P2138),
				.a2(P2148),
				.a3(P2228),
				.a4(P2238),
				.a5(P2248),
				.a6(P2328),
				.a7(P2338),
				.a8(P2348),
				.b0(W2V008),
				.b1(W2V018),
				.b2(W2V028),
				.b3(W2V108),
				.b4(W2V118),
				.b5(W2V128),
				.b6(W2V208),
				.b7(W2V218),
				.b8(W2V228),
				.c(c2812V)
);

ninexnine_unit ninexnine_unit_7517(
				.clk(clk),
				.rstn(rstn),
				.a0(P2129),
				.a1(P2139),
				.a2(P2149),
				.a3(P2229),
				.a4(P2239),
				.a5(P2249),
				.a6(P2329),
				.a7(P2339),
				.a8(P2349),
				.b0(W2V009),
				.b1(W2V019),
				.b2(W2V029),
				.b3(W2V109),
				.b4(W2V119),
				.b5(W2V129),
				.b6(W2V209),
				.b7(W2V219),
				.b8(W2V229),
				.c(c2912V)
);

ninexnine_unit ninexnine_unit_7518(
				.clk(clk),
				.rstn(rstn),
				.a0(P212A),
				.a1(P213A),
				.a2(P214A),
				.a3(P222A),
				.a4(P223A),
				.a5(P224A),
				.a6(P232A),
				.a7(P233A),
				.a8(P234A),
				.b0(W2V00A),
				.b1(W2V01A),
				.b2(W2V02A),
				.b3(W2V10A),
				.b4(W2V11A),
				.b5(W2V12A),
				.b6(W2V20A),
				.b7(W2V21A),
				.b8(W2V22A),
				.c(c2A12V)
);

ninexnine_unit ninexnine_unit_7519(
				.clk(clk),
				.rstn(rstn),
				.a0(P212B),
				.a1(P213B),
				.a2(P214B),
				.a3(P222B),
				.a4(P223B),
				.a5(P224B),
				.a6(P232B),
				.a7(P233B),
				.a8(P234B),
				.b0(W2V00B),
				.b1(W2V01B),
				.b2(W2V02B),
				.b3(W2V10B),
				.b4(W2V11B),
				.b5(W2V12B),
				.b6(W2V20B),
				.b7(W2V21B),
				.b8(W2V22B),
				.c(c2B12V)
);

ninexnine_unit ninexnine_unit_7520(
				.clk(clk),
				.rstn(rstn),
				.a0(P212C),
				.a1(P213C),
				.a2(P214C),
				.a3(P222C),
				.a4(P223C),
				.a5(P224C),
				.a6(P232C),
				.a7(P233C),
				.a8(P234C),
				.b0(W2V00C),
				.b1(W2V01C),
				.b2(W2V02C),
				.b3(W2V10C),
				.b4(W2V11C),
				.b5(W2V12C),
				.b6(W2V20C),
				.b7(W2V21C),
				.b8(W2V22C),
				.c(c2C12V)
);

ninexnine_unit ninexnine_unit_7521(
				.clk(clk),
				.rstn(rstn),
				.a0(P212D),
				.a1(P213D),
				.a2(P214D),
				.a3(P222D),
				.a4(P223D),
				.a5(P224D),
				.a6(P232D),
				.a7(P233D),
				.a8(P234D),
				.b0(W2V00D),
				.b1(W2V01D),
				.b2(W2V02D),
				.b3(W2V10D),
				.b4(W2V11D),
				.b5(W2V12D),
				.b6(W2V20D),
				.b7(W2V21D),
				.b8(W2V22D),
				.c(c2D12V)
);

ninexnine_unit ninexnine_unit_7522(
				.clk(clk),
				.rstn(rstn),
				.a0(P212E),
				.a1(P213E),
				.a2(P214E),
				.a3(P222E),
				.a4(P223E),
				.a5(P224E),
				.a6(P232E),
				.a7(P233E),
				.a8(P234E),
				.b0(W2V00E),
				.b1(W2V01E),
				.b2(W2V02E),
				.b3(W2V10E),
				.b4(W2V11E),
				.b5(W2V12E),
				.b6(W2V20E),
				.b7(W2V21E),
				.b8(W2V22E),
				.c(c2E12V)
);

ninexnine_unit ninexnine_unit_7523(
				.clk(clk),
				.rstn(rstn),
				.a0(P212F),
				.a1(P213F),
				.a2(P214F),
				.a3(P222F),
				.a4(P223F),
				.a5(P224F),
				.a6(P232F),
				.a7(P233F),
				.a8(P234F),
				.b0(W2V00F),
				.b1(W2V01F),
				.b2(W2V02F),
				.b3(W2V10F),
				.b4(W2V11F),
				.b5(W2V12F),
				.b6(W2V20F),
				.b7(W2V21F),
				.b8(W2V22F),
				.c(c2F12V)
);

assign C212V=c2012V+c2112V+c2212V+c2312V+c2412V+c2512V+c2612V+c2712V+c2812V+c2912V+c2A12V+c2B12V+c2C12V+c2D12V+c2E12V+c2F12V;
assign A212V=(C212V>=0)?1:0;

assign P312V=A212V;

ninexnine_unit ninexnine_unit_7524(
				.clk(clk),
				.rstn(rstn),
				.a0(P2200),
				.a1(P2210),
				.a2(P2220),
				.a3(P2300),
				.a4(P2310),
				.a5(P2320),
				.a6(P2400),
				.a7(P2410),
				.a8(P2420),
				.b0(W2V000),
				.b1(W2V010),
				.b2(W2V020),
				.b3(W2V100),
				.b4(W2V110),
				.b5(W2V120),
				.b6(W2V200),
				.b7(W2V210),
				.b8(W2V220),
				.c(c2020V)
);

ninexnine_unit ninexnine_unit_7525(
				.clk(clk),
				.rstn(rstn),
				.a0(P2201),
				.a1(P2211),
				.a2(P2221),
				.a3(P2301),
				.a4(P2311),
				.a5(P2321),
				.a6(P2401),
				.a7(P2411),
				.a8(P2421),
				.b0(W2V001),
				.b1(W2V011),
				.b2(W2V021),
				.b3(W2V101),
				.b4(W2V111),
				.b5(W2V121),
				.b6(W2V201),
				.b7(W2V211),
				.b8(W2V221),
				.c(c2120V)
);

ninexnine_unit ninexnine_unit_7526(
				.clk(clk),
				.rstn(rstn),
				.a0(P2202),
				.a1(P2212),
				.a2(P2222),
				.a3(P2302),
				.a4(P2312),
				.a5(P2322),
				.a6(P2402),
				.a7(P2412),
				.a8(P2422),
				.b0(W2V002),
				.b1(W2V012),
				.b2(W2V022),
				.b3(W2V102),
				.b4(W2V112),
				.b5(W2V122),
				.b6(W2V202),
				.b7(W2V212),
				.b8(W2V222),
				.c(c2220V)
);

ninexnine_unit ninexnine_unit_7527(
				.clk(clk),
				.rstn(rstn),
				.a0(P2203),
				.a1(P2213),
				.a2(P2223),
				.a3(P2303),
				.a4(P2313),
				.a5(P2323),
				.a6(P2403),
				.a7(P2413),
				.a8(P2423),
				.b0(W2V003),
				.b1(W2V013),
				.b2(W2V023),
				.b3(W2V103),
				.b4(W2V113),
				.b5(W2V123),
				.b6(W2V203),
				.b7(W2V213),
				.b8(W2V223),
				.c(c2320V)
);

ninexnine_unit ninexnine_unit_7528(
				.clk(clk),
				.rstn(rstn),
				.a0(P2204),
				.a1(P2214),
				.a2(P2224),
				.a3(P2304),
				.a4(P2314),
				.a5(P2324),
				.a6(P2404),
				.a7(P2414),
				.a8(P2424),
				.b0(W2V004),
				.b1(W2V014),
				.b2(W2V024),
				.b3(W2V104),
				.b4(W2V114),
				.b5(W2V124),
				.b6(W2V204),
				.b7(W2V214),
				.b8(W2V224),
				.c(c2420V)
);

ninexnine_unit ninexnine_unit_7529(
				.clk(clk),
				.rstn(rstn),
				.a0(P2205),
				.a1(P2215),
				.a2(P2225),
				.a3(P2305),
				.a4(P2315),
				.a5(P2325),
				.a6(P2405),
				.a7(P2415),
				.a8(P2425),
				.b0(W2V005),
				.b1(W2V015),
				.b2(W2V025),
				.b3(W2V105),
				.b4(W2V115),
				.b5(W2V125),
				.b6(W2V205),
				.b7(W2V215),
				.b8(W2V225),
				.c(c2520V)
);

ninexnine_unit ninexnine_unit_7530(
				.clk(clk),
				.rstn(rstn),
				.a0(P2206),
				.a1(P2216),
				.a2(P2226),
				.a3(P2306),
				.a4(P2316),
				.a5(P2326),
				.a6(P2406),
				.a7(P2416),
				.a8(P2426),
				.b0(W2V006),
				.b1(W2V016),
				.b2(W2V026),
				.b3(W2V106),
				.b4(W2V116),
				.b5(W2V126),
				.b6(W2V206),
				.b7(W2V216),
				.b8(W2V226),
				.c(c2620V)
);

ninexnine_unit ninexnine_unit_7531(
				.clk(clk),
				.rstn(rstn),
				.a0(P2207),
				.a1(P2217),
				.a2(P2227),
				.a3(P2307),
				.a4(P2317),
				.a5(P2327),
				.a6(P2407),
				.a7(P2417),
				.a8(P2427),
				.b0(W2V007),
				.b1(W2V017),
				.b2(W2V027),
				.b3(W2V107),
				.b4(W2V117),
				.b5(W2V127),
				.b6(W2V207),
				.b7(W2V217),
				.b8(W2V227),
				.c(c2720V)
);

ninexnine_unit ninexnine_unit_7532(
				.clk(clk),
				.rstn(rstn),
				.a0(P2208),
				.a1(P2218),
				.a2(P2228),
				.a3(P2308),
				.a4(P2318),
				.a5(P2328),
				.a6(P2408),
				.a7(P2418),
				.a8(P2428),
				.b0(W2V008),
				.b1(W2V018),
				.b2(W2V028),
				.b3(W2V108),
				.b4(W2V118),
				.b5(W2V128),
				.b6(W2V208),
				.b7(W2V218),
				.b8(W2V228),
				.c(c2820V)
);

ninexnine_unit ninexnine_unit_7533(
				.clk(clk),
				.rstn(rstn),
				.a0(P2209),
				.a1(P2219),
				.a2(P2229),
				.a3(P2309),
				.a4(P2319),
				.a5(P2329),
				.a6(P2409),
				.a7(P2419),
				.a8(P2429),
				.b0(W2V009),
				.b1(W2V019),
				.b2(W2V029),
				.b3(W2V109),
				.b4(W2V119),
				.b5(W2V129),
				.b6(W2V209),
				.b7(W2V219),
				.b8(W2V229),
				.c(c2920V)
);

ninexnine_unit ninexnine_unit_7534(
				.clk(clk),
				.rstn(rstn),
				.a0(P220A),
				.a1(P221A),
				.a2(P222A),
				.a3(P230A),
				.a4(P231A),
				.a5(P232A),
				.a6(P240A),
				.a7(P241A),
				.a8(P242A),
				.b0(W2V00A),
				.b1(W2V01A),
				.b2(W2V02A),
				.b3(W2V10A),
				.b4(W2V11A),
				.b5(W2V12A),
				.b6(W2V20A),
				.b7(W2V21A),
				.b8(W2V22A),
				.c(c2A20V)
);

ninexnine_unit ninexnine_unit_7535(
				.clk(clk),
				.rstn(rstn),
				.a0(P220B),
				.a1(P221B),
				.a2(P222B),
				.a3(P230B),
				.a4(P231B),
				.a5(P232B),
				.a6(P240B),
				.a7(P241B),
				.a8(P242B),
				.b0(W2V00B),
				.b1(W2V01B),
				.b2(W2V02B),
				.b3(W2V10B),
				.b4(W2V11B),
				.b5(W2V12B),
				.b6(W2V20B),
				.b7(W2V21B),
				.b8(W2V22B),
				.c(c2B20V)
);

ninexnine_unit ninexnine_unit_7536(
				.clk(clk),
				.rstn(rstn),
				.a0(P220C),
				.a1(P221C),
				.a2(P222C),
				.a3(P230C),
				.a4(P231C),
				.a5(P232C),
				.a6(P240C),
				.a7(P241C),
				.a8(P242C),
				.b0(W2V00C),
				.b1(W2V01C),
				.b2(W2V02C),
				.b3(W2V10C),
				.b4(W2V11C),
				.b5(W2V12C),
				.b6(W2V20C),
				.b7(W2V21C),
				.b8(W2V22C),
				.c(c2C20V)
);

ninexnine_unit ninexnine_unit_7537(
				.clk(clk),
				.rstn(rstn),
				.a0(P220D),
				.a1(P221D),
				.a2(P222D),
				.a3(P230D),
				.a4(P231D),
				.a5(P232D),
				.a6(P240D),
				.a7(P241D),
				.a8(P242D),
				.b0(W2V00D),
				.b1(W2V01D),
				.b2(W2V02D),
				.b3(W2V10D),
				.b4(W2V11D),
				.b5(W2V12D),
				.b6(W2V20D),
				.b7(W2V21D),
				.b8(W2V22D),
				.c(c2D20V)
);

ninexnine_unit ninexnine_unit_7538(
				.clk(clk),
				.rstn(rstn),
				.a0(P220E),
				.a1(P221E),
				.a2(P222E),
				.a3(P230E),
				.a4(P231E),
				.a5(P232E),
				.a6(P240E),
				.a7(P241E),
				.a8(P242E),
				.b0(W2V00E),
				.b1(W2V01E),
				.b2(W2V02E),
				.b3(W2V10E),
				.b4(W2V11E),
				.b5(W2V12E),
				.b6(W2V20E),
				.b7(W2V21E),
				.b8(W2V22E),
				.c(c2E20V)
);

ninexnine_unit ninexnine_unit_7539(
				.clk(clk),
				.rstn(rstn),
				.a0(P220F),
				.a1(P221F),
				.a2(P222F),
				.a3(P230F),
				.a4(P231F),
				.a5(P232F),
				.a6(P240F),
				.a7(P241F),
				.a8(P242F),
				.b0(W2V00F),
				.b1(W2V01F),
				.b2(W2V02F),
				.b3(W2V10F),
				.b4(W2V11F),
				.b5(W2V12F),
				.b6(W2V20F),
				.b7(W2V21F),
				.b8(W2V22F),
				.c(c2F20V)
);

assign C220V=c2020V+c2120V+c2220V+c2320V+c2420V+c2520V+c2620V+c2720V+c2820V+c2920V+c2A20V+c2B20V+c2C20V+c2D20V+c2E20V+c2F20V;
assign A220V=(C220V>=0)?1:0;

assign P320V=A220V;

ninexnine_unit ninexnine_unit_7540(
				.clk(clk),
				.rstn(rstn),
				.a0(P2210),
				.a1(P2220),
				.a2(P2230),
				.a3(P2310),
				.a4(P2320),
				.a5(P2330),
				.a6(P2410),
				.a7(P2420),
				.a8(P2430),
				.b0(W2V000),
				.b1(W2V010),
				.b2(W2V020),
				.b3(W2V100),
				.b4(W2V110),
				.b5(W2V120),
				.b6(W2V200),
				.b7(W2V210),
				.b8(W2V220),
				.c(c2021V)
);

ninexnine_unit ninexnine_unit_7541(
				.clk(clk),
				.rstn(rstn),
				.a0(P2211),
				.a1(P2221),
				.a2(P2231),
				.a3(P2311),
				.a4(P2321),
				.a5(P2331),
				.a6(P2411),
				.a7(P2421),
				.a8(P2431),
				.b0(W2V001),
				.b1(W2V011),
				.b2(W2V021),
				.b3(W2V101),
				.b4(W2V111),
				.b5(W2V121),
				.b6(W2V201),
				.b7(W2V211),
				.b8(W2V221),
				.c(c2121V)
);

ninexnine_unit ninexnine_unit_7542(
				.clk(clk),
				.rstn(rstn),
				.a0(P2212),
				.a1(P2222),
				.a2(P2232),
				.a3(P2312),
				.a4(P2322),
				.a5(P2332),
				.a6(P2412),
				.a7(P2422),
				.a8(P2432),
				.b0(W2V002),
				.b1(W2V012),
				.b2(W2V022),
				.b3(W2V102),
				.b4(W2V112),
				.b5(W2V122),
				.b6(W2V202),
				.b7(W2V212),
				.b8(W2V222),
				.c(c2221V)
);

ninexnine_unit ninexnine_unit_7543(
				.clk(clk),
				.rstn(rstn),
				.a0(P2213),
				.a1(P2223),
				.a2(P2233),
				.a3(P2313),
				.a4(P2323),
				.a5(P2333),
				.a6(P2413),
				.a7(P2423),
				.a8(P2433),
				.b0(W2V003),
				.b1(W2V013),
				.b2(W2V023),
				.b3(W2V103),
				.b4(W2V113),
				.b5(W2V123),
				.b6(W2V203),
				.b7(W2V213),
				.b8(W2V223),
				.c(c2321V)
);

ninexnine_unit ninexnine_unit_7544(
				.clk(clk),
				.rstn(rstn),
				.a0(P2214),
				.a1(P2224),
				.a2(P2234),
				.a3(P2314),
				.a4(P2324),
				.a5(P2334),
				.a6(P2414),
				.a7(P2424),
				.a8(P2434),
				.b0(W2V004),
				.b1(W2V014),
				.b2(W2V024),
				.b3(W2V104),
				.b4(W2V114),
				.b5(W2V124),
				.b6(W2V204),
				.b7(W2V214),
				.b8(W2V224),
				.c(c2421V)
);

ninexnine_unit ninexnine_unit_7545(
				.clk(clk),
				.rstn(rstn),
				.a0(P2215),
				.a1(P2225),
				.a2(P2235),
				.a3(P2315),
				.a4(P2325),
				.a5(P2335),
				.a6(P2415),
				.a7(P2425),
				.a8(P2435),
				.b0(W2V005),
				.b1(W2V015),
				.b2(W2V025),
				.b3(W2V105),
				.b4(W2V115),
				.b5(W2V125),
				.b6(W2V205),
				.b7(W2V215),
				.b8(W2V225),
				.c(c2521V)
);

ninexnine_unit ninexnine_unit_7546(
				.clk(clk),
				.rstn(rstn),
				.a0(P2216),
				.a1(P2226),
				.a2(P2236),
				.a3(P2316),
				.a4(P2326),
				.a5(P2336),
				.a6(P2416),
				.a7(P2426),
				.a8(P2436),
				.b0(W2V006),
				.b1(W2V016),
				.b2(W2V026),
				.b3(W2V106),
				.b4(W2V116),
				.b5(W2V126),
				.b6(W2V206),
				.b7(W2V216),
				.b8(W2V226),
				.c(c2621V)
);

ninexnine_unit ninexnine_unit_7547(
				.clk(clk),
				.rstn(rstn),
				.a0(P2217),
				.a1(P2227),
				.a2(P2237),
				.a3(P2317),
				.a4(P2327),
				.a5(P2337),
				.a6(P2417),
				.a7(P2427),
				.a8(P2437),
				.b0(W2V007),
				.b1(W2V017),
				.b2(W2V027),
				.b3(W2V107),
				.b4(W2V117),
				.b5(W2V127),
				.b6(W2V207),
				.b7(W2V217),
				.b8(W2V227),
				.c(c2721V)
);

ninexnine_unit ninexnine_unit_7548(
				.clk(clk),
				.rstn(rstn),
				.a0(P2218),
				.a1(P2228),
				.a2(P2238),
				.a3(P2318),
				.a4(P2328),
				.a5(P2338),
				.a6(P2418),
				.a7(P2428),
				.a8(P2438),
				.b0(W2V008),
				.b1(W2V018),
				.b2(W2V028),
				.b3(W2V108),
				.b4(W2V118),
				.b5(W2V128),
				.b6(W2V208),
				.b7(W2V218),
				.b8(W2V228),
				.c(c2821V)
);

ninexnine_unit ninexnine_unit_7549(
				.clk(clk),
				.rstn(rstn),
				.a0(P2219),
				.a1(P2229),
				.a2(P2239),
				.a3(P2319),
				.a4(P2329),
				.a5(P2339),
				.a6(P2419),
				.a7(P2429),
				.a8(P2439),
				.b0(W2V009),
				.b1(W2V019),
				.b2(W2V029),
				.b3(W2V109),
				.b4(W2V119),
				.b5(W2V129),
				.b6(W2V209),
				.b7(W2V219),
				.b8(W2V229),
				.c(c2921V)
);

ninexnine_unit ninexnine_unit_7550(
				.clk(clk),
				.rstn(rstn),
				.a0(P221A),
				.a1(P222A),
				.a2(P223A),
				.a3(P231A),
				.a4(P232A),
				.a5(P233A),
				.a6(P241A),
				.a7(P242A),
				.a8(P243A),
				.b0(W2V00A),
				.b1(W2V01A),
				.b2(W2V02A),
				.b3(W2V10A),
				.b4(W2V11A),
				.b5(W2V12A),
				.b6(W2V20A),
				.b7(W2V21A),
				.b8(W2V22A),
				.c(c2A21V)
);

ninexnine_unit ninexnine_unit_7551(
				.clk(clk),
				.rstn(rstn),
				.a0(P221B),
				.a1(P222B),
				.a2(P223B),
				.a3(P231B),
				.a4(P232B),
				.a5(P233B),
				.a6(P241B),
				.a7(P242B),
				.a8(P243B),
				.b0(W2V00B),
				.b1(W2V01B),
				.b2(W2V02B),
				.b3(W2V10B),
				.b4(W2V11B),
				.b5(W2V12B),
				.b6(W2V20B),
				.b7(W2V21B),
				.b8(W2V22B),
				.c(c2B21V)
);

ninexnine_unit ninexnine_unit_7552(
				.clk(clk),
				.rstn(rstn),
				.a0(P221C),
				.a1(P222C),
				.a2(P223C),
				.a3(P231C),
				.a4(P232C),
				.a5(P233C),
				.a6(P241C),
				.a7(P242C),
				.a8(P243C),
				.b0(W2V00C),
				.b1(W2V01C),
				.b2(W2V02C),
				.b3(W2V10C),
				.b4(W2V11C),
				.b5(W2V12C),
				.b6(W2V20C),
				.b7(W2V21C),
				.b8(W2V22C),
				.c(c2C21V)
);

ninexnine_unit ninexnine_unit_7553(
				.clk(clk),
				.rstn(rstn),
				.a0(P221D),
				.a1(P222D),
				.a2(P223D),
				.a3(P231D),
				.a4(P232D),
				.a5(P233D),
				.a6(P241D),
				.a7(P242D),
				.a8(P243D),
				.b0(W2V00D),
				.b1(W2V01D),
				.b2(W2V02D),
				.b3(W2V10D),
				.b4(W2V11D),
				.b5(W2V12D),
				.b6(W2V20D),
				.b7(W2V21D),
				.b8(W2V22D),
				.c(c2D21V)
);

ninexnine_unit ninexnine_unit_7554(
				.clk(clk),
				.rstn(rstn),
				.a0(P221E),
				.a1(P222E),
				.a2(P223E),
				.a3(P231E),
				.a4(P232E),
				.a5(P233E),
				.a6(P241E),
				.a7(P242E),
				.a8(P243E),
				.b0(W2V00E),
				.b1(W2V01E),
				.b2(W2V02E),
				.b3(W2V10E),
				.b4(W2V11E),
				.b5(W2V12E),
				.b6(W2V20E),
				.b7(W2V21E),
				.b8(W2V22E),
				.c(c2E21V)
);

ninexnine_unit ninexnine_unit_7555(
				.clk(clk),
				.rstn(rstn),
				.a0(P221F),
				.a1(P222F),
				.a2(P223F),
				.a3(P231F),
				.a4(P232F),
				.a5(P233F),
				.a6(P241F),
				.a7(P242F),
				.a8(P243F),
				.b0(W2V00F),
				.b1(W2V01F),
				.b2(W2V02F),
				.b3(W2V10F),
				.b4(W2V11F),
				.b5(W2V12F),
				.b6(W2V20F),
				.b7(W2V21F),
				.b8(W2V22F),
				.c(c2F21V)
);

assign C221V=c2021V+c2121V+c2221V+c2321V+c2421V+c2521V+c2621V+c2721V+c2821V+c2921V+c2A21V+c2B21V+c2C21V+c2D21V+c2E21V+c2F21V;
assign A221V=(C221V>=0)?1:0;

assign P321V=A221V;

ninexnine_unit ninexnine_unit_7556(
				.clk(clk),
				.rstn(rstn),
				.a0(P2220),
				.a1(P2230),
				.a2(P2240),
				.a3(P2320),
				.a4(P2330),
				.a5(P2340),
				.a6(P2420),
				.a7(P2430),
				.a8(P2440),
				.b0(W2V000),
				.b1(W2V010),
				.b2(W2V020),
				.b3(W2V100),
				.b4(W2V110),
				.b5(W2V120),
				.b6(W2V200),
				.b7(W2V210),
				.b8(W2V220),
				.c(c2022V)
);

ninexnine_unit ninexnine_unit_7557(
				.clk(clk),
				.rstn(rstn),
				.a0(P2221),
				.a1(P2231),
				.a2(P2241),
				.a3(P2321),
				.a4(P2331),
				.a5(P2341),
				.a6(P2421),
				.a7(P2431),
				.a8(P2441),
				.b0(W2V001),
				.b1(W2V011),
				.b2(W2V021),
				.b3(W2V101),
				.b4(W2V111),
				.b5(W2V121),
				.b6(W2V201),
				.b7(W2V211),
				.b8(W2V221),
				.c(c2122V)
);

ninexnine_unit ninexnine_unit_7558(
				.clk(clk),
				.rstn(rstn),
				.a0(P2222),
				.a1(P2232),
				.a2(P2242),
				.a3(P2322),
				.a4(P2332),
				.a5(P2342),
				.a6(P2422),
				.a7(P2432),
				.a8(P2442),
				.b0(W2V002),
				.b1(W2V012),
				.b2(W2V022),
				.b3(W2V102),
				.b4(W2V112),
				.b5(W2V122),
				.b6(W2V202),
				.b7(W2V212),
				.b8(W2V222),
				.c(c2222V)
);

ninexnine_unit ninexnine_unit_7559(
				.clk(clk),
				.rstn(rstn),
				.a0(P2223),
				.a1(P2233),
				.a2(P2243),
				.a3(P2323),
				.a4(P2333),
				.a5(P2343),
				.a6(P2423),
				.a7(P2433),
				.a8(P2443),
				.b0(W2V003),
				.b1(W2V013),
				.b2(W2V023),
				.b3(W2V103),
				.b4(W2V113),
				.b5(W2V123),
				.b6(W2V203),
				.b7(W2V213),
				.b8(W2V223),
				.c(c2322V)
);

ninexnine_unit ninexnine_unit_7560(
				.clk(clk),
				.rstn(rstn),
				.a0(P2224),
				.a1(P2234),
				.a2(P2244),
				.a3(P2324),
				.a4(P2334),
				.a5(P2344),
				.a6(P2424),
				.a7(P2434),
				.a8(P2444),
				.b0(W2V004),
				.b1(W2V014),
				.b2(W2V024),
				.b3(W2V104),
				.b4(W2V114),
				.b5(W2V124),
				.b6(W2V204),
				.b7(W2V214),
				.b8(W2V224),
				.c(c2422V)
);

ninexnine_unit ninexnine_unit_7561(
				.clk(clk),
				.rstn(rstn),
				.a0(P2225),
				.a1(P2235),
				.a2(P2245),
				.a3(P2325),
				.a4(P2335),
				.a5(P2345),
				.a6(P2425),
				.a7(P2435),
				.a8(P2445),
				.b0(W2V005),
				.b1(W2V015),
				.b2(W2V025),
				.b3(W2V105),
				.b4(W2V115),
				.b5(W2V125),
				.b6(W2V205),
				.b7(W2V215),
				.b8(W2V225),
				.c(c2522V)
);

ninexnine_unit ninexnine_unit_7562(
				.clk(clk),
				.rstn(rstn),
				.a0(P2226),
				.a1(P2236),
				.a2(P2246),
				.a3(P2326),
				.a4(P2336),
				.a5(P2346),
				.a6(P2426),
				.a7(P2436),
				.a8(P2446),
				.b0(W2V006),
				.b1(W2V016),
				.b2(W2V026),
				.b3(W2V106),
				.b4(W2V116),
				.b5(W2V126),
				.b6(W2V206),
				.b7(W2V216),
				.b8(W2V226),
				.c(c2622V)
);

ninexnine_unit ninexnine_unit_7563(
				.clk(clk),
				.rstn(rstn),
				.a0(P2227),
				.a1(P2237),
				.a2(P2247),
				.a3(P2327),
				.a4(P2337),
				.a5(P2347),
				.a6(P2427),
				.a7(P2437),
				.a8(P2447),
				.b0(W2V007),
				.b1(W2V017),
				.b2(W2V027),
				.b3(W2V107),
				.b4(W2V117),
				.b5(W2V127),
				.b6(W2V207),
				.b7(W2V217),
				.b8(W2V227),
				.c(c2722V)
);

ninexnine_unit ninexnine_unit_7564(
				.clk(clk),
				.rstn(rstn),
				.a0(P2228),
				.a1(P2238),
				.a2(P2248),
				.a3(P2328),
				.a4(P2338),
				.a5(P2348),
				.a6(P2428),
				.a7(P2438),
				.a8(P2448),
				.b0(W2V008),
				.b1(W2V018),
				.b2(W2V028),
				.b3(W2V108),
				.b4(W2V118),
				.b5(W2V128),
				.b6(W2V208),
				.b7(W2V218),
				.b8(W2V228),
				.c(c2822V)
);

ninexnine_unit ninexnine_unit_7565(
				.clk(clk),
				.rstn(rstn),
				.a0(P2229),
				.a1(P2239),
				.a2(P2249),
				.a3(P2329),
				.a4(P2339),
				.a5(P2349),
				.a6(P2429),
				.a7(P2439),
				.a8(P2449),
				.b0(W2V009),
				.b1(W2V019),
				.b2(W2V029),
				.b3(W2V109),
				.b4(W2V119),
				.b5(W2V129),
				.b6(W2V209),
				.b7(W2V219),
				.b8(W2V229),
				.c(c2922V)
);

ninexnine_unit ninexnine_unit_7566(
				.clk(clk),
				.rstn(rstn),
				.a0(P222A),
				.a1(P223A),
				.a2(P224A),
				.a3(P232A),
				.a4(P233A),
				.a5(P234A),
				.a6(P242A),
				.a7(P243A),
				.a8(P244A),
				.b0(W2V00A),
				.b1(W2V01A),
				.b2(W2V02A),
				.b3(W2V10A),
				.b4(W2V11A),
				.b5(W2V12A),
				.b6(W2V20A),
				.b7(W2V21A),
				.b8(W2V22A),
				.c(c2A22V)
);

ninexnine_unit ninexnine_unit_7567(
				.clk(clk),
				.rstn(rstn),
				.a0(P222B),
				.a1(P223B),
				.a2(P224B),
				.a3(P232B),
				.a4(P233B),
				.a5(P234B),
				.a6(P242B),
				.a7(P243B),
				.a8(P244B),
				.b0(W2V00B),
				.b1(W2V01B),
				.b2(W2V02B),
				.b3(W2V10B),
				.b4(W2V11B),
				.b5(W2V12B),
				.b6(W2V20B),
				.b7(W2V21B),
				.b8(W2V22B),
				.c(c2B22V)
);

ninexnine_unit ninexnine_unit_7568(
				.clk(clk),
				.rstn(rstn),
				.a0(P222C),
				.a1(P223C),
				.a2(P224C),
				.a3(P232C),
				.a4(P233C),
				.a5(P234C),
				.a6(P242C),
				.a7(P243C),
				.a8(P244C),
				.b0(W2V00C),
				.b1(W2V01C),
				.b2(W2V02C),
				.b3(W2V10C),
				.b4(W2V11C),
				.b5(W2V12C),
				.b6(W2V20C),
				.b7(W2V21C),
				.b8(W2V22C),
				.c(c2C22V)
);

ninexnine_unit ninexnine_unit_7569(
				.clk(clk),
				.rstn(rstn),
				.a0(P222D),
				.a1(P223D),
				.a2(P224D),
				.a3(P232D),
				.a4(P233D),
				.a5(P234D),
				.a6(P242D),
				.a7(P243D),
				.a8(P244D),
				.b0(W2V00D),
				.b1(W2V01D),
				.b2(W2V02D),
				.b3(W2V10D),
				.b4(W2V11D),
				.b5(W2V12D),
				.b6(W2V20D),
				.b7(W2V21D),
				.b8(W2V22D),
				.c(c2D22V)
);

ninexnine_unit ninexnine_unit_7570(
				.clk(clk),
				.rstn(rstn),
				.a0(P222E),
				.a1(P223E),
				.a2(P224E),
				.a3(P232E),
				.a4(P233E),
				.a5(P234E),
				.a6(P242E),
				.a7(P243E),
				.a8(P244E),
				.b0(W2V00E),
				.b1(W2V01E),
				.b2(W2V02E),
				.b3(W2V10E),
				.b4(W2V11E),
				.b5(W2V12E),
				.b6(W2V20E),
				.b7(W2V21E),
				.b8(W2V22E),
				.c(c2E22V)
);

ninexnine_unit ninexnine_unit_7571(
				.clk(clk),
				.rstn(rstn),
				.a0(P222F),
				.a1(P223F),
				.a2(P224F),
				.a3(P232F),
				.a4(P233F),
				.a5(P234F),
				.a6(P242F),
				.a7(P243F),
				.a8(P244F),
				.b0(W2V00F),
				.b1(W2V01F),
				.b2(W2V02F),
				.b3(W2V10F),
				.b4(W2V11F),
				.b5(W2V12F),
				.b6(W2V20F),
				.b7(W2V21F),
				.b8(W2V22F),
				.c(c2F22V)
);

assign C222V=c2022V+c2122V+c2222V+c2322V+c2422V+c2522V+c2622V+c2722V+c2822V+c2922V+c2A22V+c2B22V+c2C22V+c2D22V+c2E22V+c2F22V;
assign A222V=(C222V>=0)?1:0;

assign P322V=A222V;

//layer3 done, begain next layer
wire P4000;
wire P4001;
wire W30000,W30010,W30020,W30100,W30110,W30120,W30200,W30210,W30220;
wire W30001,W30011,W30021,W30101,W30111,W30121,W30201,W30211,W30221;
wire W30002,W30012,W30022,W30102,W30112,W30122,W30202,W30212,W30222;
wire W30003,W30013,W30023,W30103,W30113,W30123,W30203,W30213,W30223;
wire W30004,W30014,W30024,W30104,W30114,W30124,W30204,W30214,W30224;
wire W30005,W30015,W30025,W30105,W30115,W30125,W30205,W30215,W30225;
wire W30006,W30016,W30026,W30106,W30116,W30126,W30206,W30216,W30226;
wire W30007,W30017,W30027,W30107,W30117,W30127,W30207,W30217,W30227;
wire W30008,W30018,W30028,W30108,W30118,W30128,W30208,W30218,W30228;
wire W30009,W30019,W30029,W30109,W30119,W30129,W30209,W30219,W30229;
wire W3000A,W3001A,W3002A,W3010A,W3011A,W3012A,W3020A,W3021A,W3022A;
wire W3000B,W3001B,W3002B,W3010B,W3011B,W3012B,W3020B,W3021B,W3022B;
wire W3000C,W3001C,W3002C,W3010C,W3011C,W3012C,W3020C,W3021C,W3022C;
wire W3000D,W3001D,W3002D,W3010D,W3011D,W3012D,W3020D,W3021D,W3022D;
wire W3000E,W3001E,W3002E,W3010E,W3011E,W3012E,W3020E,W3021E,W3022E;
wire W3000F,W3001F,W3002F,W3010F,W3011F,W3012F,W3020F,W3021F,W3022F;
wire W3000G,W3001G,W3002G,W3010G,W3011G,W3012G,W3020G,W3021G,W3022G;
wire W3000H,W3001H,W3002H,W3010H,W3011H,W3012H,W3020H,W3021H,W3022H;
wire W3000I,W3001I,W3002I,W3010I,W3011I,W3012I,W3020I,W3021I,W3022I;
wire W3000J,W3001J,W3002J,W3010J,W3011J,W3012J,W3020J,W3021J,W3022J;
wire W3000K,W3001K,W3002K,W3010K,W3011K,W3012K,W3020K,W3021K,W3022K;
wire W3000L,W3001L,W3002L,W3010L,W3011L,W3012L,W3020L,W3021L,W3022L;
wire W3000M,W3001M,W3002M,W3010M,W3011M,W3012M,W3020M,W3021M,W3022M;
wire W3000N,W3001N,W3002N,W3010N,W3011N,W3012N,W3020N,W3021N,W3022N;
wire W3000O,W3001O,W3002O,W3010O,W3011O,W3012O,W3020O,W3021O,W3022O;
wire W3000P,W3001P,W3002P,W3010P,W3011P,W3012P,W3020P,W3021P,W3022P;
wire W3000Q,W3001Q,W3002Q,W3010Q,W3011Q,W3012Q,W3020Q,W3021Q,W3022Q;
wire W3000R,W3001R,W3002R,W3010R,W3011R,W3012R,W3020R,W3021R,W3022R;
wire W3000S,W3001S,W3002S,W3010S,W3011S,W3012S,W3020S,W3021S,W3022S;
wire W3000T,W3001T,W3002T,W3010T,W3011T,W3012T,W3020T,W3021T,W3022T;
wire W3000U,W3001U,W3002U,W3010U,W3011U,W3012U,W3020U,W3021U,W3022U;
wire W3000V,W3001V,W3002V,W3010V,W3011V,W3012V,W3020V,W3021V,W3022V;
wire W31000,W31010,W31020,W31100,W31110,W31120,W31200,W31210,W31220;
wire W31001,W31011,W31021,W31101,W31111,W31121,W31201,W31211,W31221;
wire W31002,W31012,W31022,W31102,W31112,W31122,W31202,W31212,W31222;
wire W31003,W31013,W31023,W31103,W31113,W31123,W31203,W31213,W31223;
wire W31004,W31014,W31024,W31104,W31114,W31124,W31204,W31214,W31224;
wire W31005,W31015,W31025,W31105,W31115,W31125,W31205,W31215,W31225;
wire W31006,W31016,W31026,W31106,W31116,W31126,W31206,W31216,W31226;
wire W31007,W31017,W31027,W31107,W31117,W31127,W31207,W31217,W31227;
wire W31008,W31018,W31028,W31108,W31118,W31128,W31208,W31218,W31228;
wire W31009,W31019,W31029,W31109,W31119,W31129,W31209,W31219,W31229;
wire W3100A,W3101A,W3102A,W3110A,W3111A,W3112A,W3120A,W3121A,W3122A;
wire W3100B,W3101B,W3102B,W3110B,W3111B,W3112B,W3120B,W3121B,W3122B;
wire W3100C,W3101C,W3102C,W3110C,W3111C,W3112C,W3120C,W3121C,W3122C;
wire W3100D,W3101D,W3102D,W3110D,W3111D,W3112D,W3120D,W3121D,W3122D;
wire W3100E,W3101E,W3102E,W3110E,W3111E,W3112E,W3120E,W3121E,W3122E;
wire W3100F,W3101F,W3102F,W3110F,W3111F,W3112F,W3120F,W3121F,W3122F;
wire W3100G,W3101G,W3102G,W3110G,W3111G,W3112G,W3120G,W3121G,W3122G;
wire W3100H,W3101H,W3102H,W3110H,W3111H,W3112H,W3120H,W3121H,W3122H;
wire W3100I,W3101I,W3102I,W3110I,W3111I,W3112I,W3120I,W3121I,W3122I;
wire W3100J,W3101J,W3102J,W3110J,W3111J,W3112J,W3120J,W3121J,W3122J;
wire W3100K,W3101K,W3102K,W3110K,W3111K,W3112K,W3120K,W3121K,W3122K;
wire W3100L,W3101L,W3102L,W3110L,W3111L,W3112L,W3120L,W3121L,W3122L;
wire W3100M,W3101M,W3102M,W3110M,W3111M,W3112M,W3120M,W3121M,W3122M;
wire W3100N,W3101N,W3102N,W3110N,W3111N,W3112N,W3120N,W3121N,W3122N;
wire W3100O,W3101O,W3102O,W3110O,W3111O,W3112O,W3120O,W3121O,W3122O;
wire W3100P,W3101P,W3102P,W3110P,W3111P,W3112P,W3120P,W3121P,W3122P;
wire W3100Q,W3101Q,W3102Q,W3110Q,W3111Q,W3112Q,W3120Q,W3121Q,W3122Q;
wire W3100R,W3101R,W3102R,W3110R,W3111R,W3112R,W3120R,W3121R,W3122R;
wire W3100S,W3101S,W3102S,W3110S,W3111S,W3112S,W3120S,W3121S,W3122S;
wire W3100T,W3101T,W3102T,W3110T,W3111T,W3112T,W3120T,W3121T,W3122T;
wire W3100U,W3101U,W3102U,W3110U,W3111U,W3112U,W3120U,W3121U,W3122U;
wire W3100V,W3101V,W3102V,W3110V,W3111V,W3112V,W3120V,W3121V,W3122V;
wire signed [4:0] c30000,c31000,c32000,c33000,c34000,c35000,c36000,c37000,c38000,c39000,c3A000,c3B000,c3C000,c3D000,c3E000,c3F000,c3G000,c3H000,c3I000,c3J000,c3K000,c3L000,c3M000,c3N000,c3O000,c3P000,c3Q000,c3R000,c3S000,c3T000,c3U000,c3V000;
wire signed [4:0] c30001,c31001,c32001,c33001,c34001,c35001,c36001,c37001,c38001,c39001,c3A001,c3B001,c3C001,c3D001,c3E001,c3F001,c3G001,c3H001,c3I001,c3J001,c3K001,c3L001,c3M001,c3N001,c3O001,c3P001,c3Q001,c3R001,c3S001,c3T001,c3U001,c3V001;
wire signed [9:0] C3000;
wire A3000;
wire signed [9:0] C3001;
wire A3001;
DFF_save_fm DFF_W5121(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30000));
DFF_save_fm DFF_W5122(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30010));
DFF_save_fm DFF_W5123(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30020));
DFF_save_fm DFF_W5124(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30100));
DFF_save_fm DFF_W5125(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30110));
DFF_save_fm DFF_W5126(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30120));
DFF_save_fm DFF_W5127(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30200));
DFF_save_fm DFF_W5128(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30210));
DFF_save_fm DFF_W5129(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30220));
DFF_save_fm DFF_W5130(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30001));
DFF_save_fm DFF_W5131(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30011));
DFF_save_fm DFF_W5132(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30021));
DFF_save_fm DFF_W5133(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30101));
DFF_save_fm DFF_W5134(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30111));
DFF_save_fm DFF_W5135(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30121));
DFF_save_fm DFF_W5136(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30201));
DFF_save_fm DFF_W5137(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30211));
DFF_save_fm DFF_W5138(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30221));
DFF_save_fm DFF_W5139(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30002));
DFF_save_fm DFF_W5140(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30012));
DFF_save_fm DFF_W5141(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30022));
DFF_save_fm DFF_W5142(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30102));
DFF_save_fm DFF_W5143(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30112));
DFF_save_fm DFF_W5144(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30122));
DFF_save_fm DFF_W5145(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30202));
DFF_save_fm DFF_W5146(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30212));
DFF_save_fm DFF_W5147(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30222));
DFF_save_fm DFF_W5148(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30003));
DFF_save_fm DFF_W5149(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30013));
DFF_save_fm DFF_W5150(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30023));
DFF_save_fm DFF_W5151(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30103));
DFF_save_fm DFF_W5152(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30113));
DFF_save_fm DFF_W5153(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30123));
DFF_save_fm DFF_W5154(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30203));
DFF_save_fm DFF_W5155(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30213));
DFF_save_fm DFF_W5156(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30223));
DFF_save_fm DFF_W5157(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30004));
DFF_save_fm DFF_W5158(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30014));
DFF_save_fm DFF_W5159(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30024));
DFF_save_fm DFF_W5160(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30104));
DFF_save_fm DFF_W5161(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30114));
DFF_save_fm DFF_W5162(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30124));
DFF_save_fm DFF_W5163(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30204));
DFF_save_fm DFF_W5164(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30214));
DFF_save_fm DFF_W5165(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30224));
DFF_save_fm DFF_W5166(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30005));
DFF_save_fm DFF_W5167(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30015));
DFF_save_fm DFF_W5168(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30025));
DFF_save_fm DFF_W5169(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30105));
DFF_save_fm DFF_W5170(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30115));
DFF_save_fm DFF_W5171(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30125));
DFF_save_fm DFF_W5172(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30205));
DFF_save_fm DFF_W5173(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30215));
DFF_save_fm DFF_W5174(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30225));
DFF_save_fm DFF_W5175(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30006));
DFF_save_fm DFF_W5176(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30016));
DFF_save_fm DFF_W5177(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30026));
DFF_save_fm DFF_W5178(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30106));
DFF_save_fm DFF_W5179(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30116));
DFF_save_fm DFF_W5180(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30126));
DFF_save_fm DFF_W5181(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30206));
DFF_save_fm DFF_W5182(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30216));
DFF_save_fm DFF_W5183(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30226));
DFF_save_fm DFF_W5184(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30007));
DFF_save_fm DFF_W5185(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30017));
DFF_save_fm DFF_W5186(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30027));
DFF_save_fm DFF_W5187(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30107));
DFF_save_fm DFF_W5188(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30117));
DFF_save_fm DFF_W5189(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30127));
DFF_save_fm DFF_W5190(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30207));
DFF_save_fm DFF_W5191(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30217));
DFF_save_fm DFF_W5192(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30227));
DFF_save_fm DFF_W5193(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30008));
DFF_save_fm DFF_W5194(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30018));
DFF_save_fm DFF_W5195(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30028));
DFF_save_fm DFF_W5196(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30108));
DFF_save_fm DFF_W5197(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30118));
DFF_save_fm DFF_W5198(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30128));
DFF_save_fm DFF_W5199(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30208));
DFF_save_fm DFF_W5200(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30218));
DFF_save_fm DFF_W5201(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30228));
DFF_save_fm DFF_W5202(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30009));
DFF_save_fm DFF_W5203(.clk(clk),.rstn(rstn),.reset_value(0),.q(W30019));
DFF_save_fm DFF_W5204(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30029));
DFF_save_fm DFF_W5205(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30109));
DFF_save_fm DFF_W5206(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30119));
DFF_save_fm DFF_W5207(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30129));
DFF_save_fm DFF_W5208(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30209));
DFF_save_fm DFF_W5209(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30219));
DFF_save_fm DFF_W5210(.clk(clk),.rstn(rstn),.reset_value(1),.q(W30229));
DFF_save_fm DFF_W5211(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3000A));
DFF_save_fm DFF_W5212(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3001A));
DFF_save_fm DFF_W5213(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3002A));
DFF_save_fm DFF_W5214(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3010A));
DFF_save_fm DFF_W5215(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3011A));
DFF_save_fm DFF_W5216(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3012A));
DFF_save_fm DFF_W5217(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3020A));
DFF_save_fm DFF_W5218(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3021A));
DFF_save_fm DFF_W5219(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3022A));
DFF_save_fm DFF_W5220(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3000B));
DFF_save_fm DFF_W5221(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3001B));
DFF_save_fm DFF_W5222(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3002B));
DFF_save_fm DFF_W5223(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3010B));
DFF_save_fm DFF_W5224(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3011B));
DFF_save_fm DFF_W5225(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3012B));
DFF_save_fm DFF_W5226(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3020B));
DFF_save_fm DFF_W5227(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3021B));
DFF_save_fm DFF_W5228(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3022B));
DFF_save_fm DFF_W5229(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3000C));
DFF_save_fm DFF_W5230(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3001C));
DFF_save_fm DFF_W5231(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3002C));
DFF_save_fm DFF_W5232(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3010C));
DFF_save_fm DFF_W5233(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3011C));
DFF_save_fm DFF_W5234(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3012C));
DFF_save_fm DFF_W5235(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3020C));
DFF_save_fm DFF_W5236(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3021C));
DFF_save_fm DFF_W5237(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3022C));
DFF_save_fm DFF_W5238(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3000D));
DFF_save_fm DFF_W5239(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3001D));
DFF_save_fm DFF_W5240(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3002D));
DFF_save_fm DFF_W5241(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3010D));
DFF_save_fm DFF_W5242(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3011D));
DFF_save_fm DFF_W5243(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3012D));
DFF_save_fm DFF_W5244(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3020D));
DFF_save_fm DFF_W5245(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3021D));
DFF_save_fm DFF_W5246(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3022D));
DFF_save_fm DFF_W5247(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3000E));
DFF_save_fm DFF_W5248(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3001E));
DFF_save_fm DFF_W5249(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3002E));
DFF_save_fm DFF_W5250(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3010E));
DFF_save_fm DFF_W5251(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3011E));
DFF_save_fm DFF_W5252(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3012E));
DFF_save_fm DFF_W5253(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3020E));
DFF_save_fm DFF_W5254(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3021E));
DFF_save_fm DFF_W5255(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3022E));
DFF_save_fm DFF_W5256(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3000F));
DFF_save_fm DFF_W5257(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3001F));
DFF_save_fm DFF_W5258(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3002F));
DFF_save_fm DFF_W5259(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3010F));
DFF_save_fm DFF_W5260(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3011F));
DFF_save_fm DFF_W5261(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3012F));
DFF_save_fm DFF_W5262(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3020F));
DFF_save_fm DFF_W5263(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3021F));
DFF_save_fm DFF_W5264(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3022F));
DFF_save_fm DFF_W5265(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3000G));
DFF_save_fm DFF_W5266(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3001G));
DFF_save_fm DFF_W5267(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3002G));
DFF_save_fm DFF_W5268(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3010G));
DFF_save_fm DFF_W5269(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3011G));
DFF_save_fm DFF_W5270(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3012G));
DFF_save_fm DFF_W5271(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3020G));
DFF_save_fm DFF_W5272(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3021G));
DFF_save_fm DFF_W5273(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3022G));
DFF_save_fm DFF_W5274(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3000H));
DFF_save_fm DFF_W5275(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3001H));
DFF_save_fm DFF_W5276(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3002H));
DFF_save_fm DFF_W5277(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3010H));
DFF_save_fm DFF_W5278(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3011H));
DFF_save_fm DFF_W5279(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3012H));
DFF_save_fm DFF_W5280(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3020H));
DFF_save_fm DFF_W5281(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3021H));
DFF_save_fm DFF_W5282(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3022H));
DFF_save_fm DFF_W5283(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3000I));
DFF_save_fm DFF_W5284(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3001I));
DFF_save_fm DFF_W5285(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3002I));
DFF_save_fm DFF_W5286(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3010I));
DFF_save_fm DFF_W5287(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3011I));
DFF_save_fm DFF_W5288(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3012I));
DFF_save_fm DFF_W5289(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3020I));
DFF_save_fm DFF_W5290(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3021I));
DFF_save_fm DFF_W5291(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3022I));
DFF_save_fm DFF_W5292(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3000J));
DFF_save_fm DFF_W5293(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3001J));
DFF_save_fm DFF_W5294(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3002J));
DFF_save_fm DFF_W5295(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3010J));
DFF_save_fm DFF_W5296(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3011J));
DFF_save_fm DFF_W5297(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3012J));
DFF_save_fm DFF_W5298(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3020J));
DFF_save_fm DFF_W5299(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3021J));
DFF_save_fm DFF_W5300(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3022J));
DFF_save_fm DFF_W5301(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3000K));
DFF_save_fm DFF_W5302(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3001K));
DFF_save_fm DFF_W5303(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3002K));
DFF_save_fm DFF_W5304(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3010K));
DFF_save_fm DFF_W5305(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3011K));
DFF_save_fm DFF_W5306(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3012K));
DFF_save_fm DFF_W5307(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3020K));
DFF_save_fm DFF_W5308(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3021K));
DFF_save_fm DFF_W5309(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3022K));
DFF_save_fm DFF_W5310(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3000L));
DFF_save_fm DFF_W5311(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3001L));
DFF_save_fm DFF_W5312(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3002L));
DFF_save_fm DFF_W5313(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3010L));
DFF_save_fm DFF_W5314(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3011L));
DFF_save_fm DFF_W5315(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3012L));
DFF_save_fm DFF_W5316(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3020L));
DFF_save_fm DFF_W5317(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3021L));
DFF_save_fm DFF_W5318(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3022L));
DFF_save_fm DFF_W5319(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3000M));
DFF_save_fm DFF_W5320(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3001M));
DFF_save_fm DFF_W5321(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3002M));
DFF_save_fm DFF_W5322(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3010M));
DFF_save_fm DFF_W5323(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3011M));
DFF_save_fm DFF_W5324(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3012M));
DFF_save_fm DFF_W5325(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3020M));
DFF_save_fm DFF_W5326(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3021M));
DFF_save_fm DFF_W5327(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3022M));
DFF_save_fm DFF_W5328(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3000N));
DFF_save_fm DFF_W5329(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3001N));
DFF_save_fm DFF_W5330(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3002N));
DFF_save_fm DFF_W5331(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3010N));
DFF_save_fm DFF_W5332(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3011N));
DFF_save_fm DFF_W5333(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3012N));
DFF_save_fm DFF_W5334(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3020N));
DFF_save_fm DFF_W5335(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3021N));
DFF_save_fm DFF_W5336(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3022N));
DFF_save_fm DFF_W5337(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3000O));
DFF_save_fm DFF_W5338(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3001O));
DFF_save_fm DFF_W5339(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3002O));
DFF_save_fm DFF_W5340(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3010O));
DFF_save_fm DFF_W5341(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3011O));
DFF_save_fm DFF_W5342(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3012O));
DFF_save_fm DFF_W5343(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3020O));
DFF_save_fm DFF_W5344(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3021O));
DFF_save_fm DFF_W5345(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3022O));
DFF_save_fm DFF_W5346(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3000P));
DFF_save_fm DFF_W5347(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3001P));
DFF_save_fm DFF_W5348(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3002P));
DFF_save_fm DFF_W5349(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3010P));
DFF_save_fm DFF_W5350(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3011P));
DFF_save_fm DFF_W5351(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3012P));
DFF_save_fm DFF_W5352(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3020P));
DFF_save_fm DFF_W5353(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3021P));
DFF_save_fm DFF_W5354(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3022P));
DFF_save_fm DFF_W5355(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3000Q));
DFF_save_fm DFF_W5356(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3001Q));
DFF_save_fm DFF_W5357(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3002Q));
DFF_save_fm DFF_W5358(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3010Q));
DFF_save_fm DFF_W5359(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3011Q));
DFF_save_fm DFF_W5360(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3012Q));
DFF_save_fm DFF_W5361(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3020Q));
DFF_save_fm DFF_W5362(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3021Q));
DFF_save_fm DFF_W5363(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3022Q));
DFF_save_fm DFF_W5364(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3000R));
DFF_save_fm DFF_W5365(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3001R));
DFF_save_fm DFF_W5366(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3002R));
DFF_save_fm DFF_W5367(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3010R));
DFF_save_fm DFF_W5368(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3011R));
DFF_save_fm DFF_W5369(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3012R));
DFF_save_fm DFF_W5370(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3020R));
DFF_save_fm DFF_W5371(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3021R));
DFF_save_fm DFF_W5372(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3022R));
DFF_save_fm DFF_W5373(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3000S));
DFF_save_fm DFF_W5374(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3001S));
DFF_save_fm DFF_W5375(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3002S));
DFF_save_fm DFF_W5376(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3010S));
DFF_save_fm DFF_W5377(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3011S));
DFF_save_fm DFF_W5378(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3012S));
DFF_save_fm DFF_W5379(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3020S));
DFF_save_fm DFF_W5380(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3021S));
DFF_save_fm DFF_W5381(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3022S));
DFF_save_fm DFF_W5382(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3000T));
DFF_save_fm DFF_W5383(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3001T));
DFF_save_fm DFF_W5384(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3002T));
DFF_save_fm DFF_W5385(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3010T));
DFF_save_fm DFF_W5386(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3011T));
DFF_save_fm DFF_W5387(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3012T));
DFF_save_fm DFF_W5388(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3020T));
DFF_save_fm DFF_W5389(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3021T));
DFF_save_fm DFF_W5390(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3022T));
DFF_save_fm DFF_W5391(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3000U));
DFF_save_fm DFF_W5392(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3001U));
DFF_save_fm DFF_W5393(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3002U));
DFF_save_fm DFF_W5394(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3010U));
DFF_save_fm DFF_W5395(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3011U));
DFF_save_fm DFF_W5396(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3012U));
DFF_save_fm DFF_W5397(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3020U));
DFF_save_fm DFF_W5398(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3021U));
DFF_save_fm DFF_W5399(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3022U));
DFF_save_fm DFF_W5400(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3000V));
DFF_save_fm DFF_W5401(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3001V));
DFF_save_fm DFF_W5402(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3002V));
DFF_save_fm DFF_W5403(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3010V));
DFF_save_fm DFF_W5404(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3011V));
DFF_save_fm DFF_W5405(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3012V));
DFF_save_fm DFF_W5406(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3020V));
DFF_save_fm DFF_W5407(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3021V));
DFF_save_fm DFF_W5408(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3022V));
DFF_save_fm DFF_W5409(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31000));
DFF_save_fm DFF_W5410(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31010));
DFF_save_fm DFF_W5411(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31020));
DFF_save_fm DFF_W5412(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31100));
DFF_save_fm DFF_W5413(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31110));
DFF_save_fm DFF_W5414(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31120));
DFF_save_fm DFF_W5415(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31200));
DFF_save_fm DFF_W5416(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31210));
DFF_save_fm DFF_W5417(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31220));
DFF_save_fm DFF_W5418(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31001));
DFF_save_fm DFF_W5419(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31011));
DFF_save_fm DFF_W5420(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31021));
DFF_save_fm DFF_W5421(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31101));
DFF_save_fm DFF_W5422(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31111));
DFF_save_fm DFF_W5423(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31121));
DFF_save_fm DFF_W5424(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31201));
DFF_save_fm DFF_W5425(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31211));
DFF_save_fm DFF_W5426(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31221));
DFF_save_fm DFF_W5427(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31002));
DFF_save_fm DFF_W5428(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31012));
DFF_save_fm DFF_W5429(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31022));
DFF_save_fm DFF_W5430(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31102));
DFF_save_fm DFF_W5431(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31112));
DFF_save_fm DFF_W5432(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31122));
DFF_save_fm DFF_W5433(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31202));
DFF_save_fm DFF_W5434(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31212));
DFF_save_fm DFF_W5435(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31222));
DFF_save_fm DFF_W5436(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31003));
DFF_save_fm DFF_W5437(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31013));
DFF_save_fm DFF_W5438(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31023));
DFF_save_fm DFF_W5439(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31103));
DFF_save_fm DFF_W5440(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31113));
DFF_save_fm DFF_W5441(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31123));
DFF_save_fm DFF_W5442(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31203));
DFF_save_fm DFF_W5443(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31213));
DFF_save_fm DFF_W5444(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31223));
DFF_save_fm DFF_W5445(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31004));
DFF_save_fm DFF_W5446(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31014));
DFF_save_fm DFF_W5447(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31024));
DFF_save_fm DFF_W5448(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31104));
DFF_save_fm DFF_W5449(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31114));
DFF_save_fm DFF_W5450(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31124));
DFF_save_fm DFF_W5451(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31204));
DFF_save_fm DFF_W5452(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31214));
DFF_save_fm DFF_W5453(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31224));
DFF_save_fm DFF_W5454(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31005));
DFF_save_fm DFF_W5455(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31015));
DFF_save_fm DFF_W5456(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31025));
DFF_save_fm DFF_W5457(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31105));
DFF_save_fm DFF_W5458(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31115));
DFF_save_fm DFF_W5459(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31125));
DFF_save_fm DFF_W5460(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31205));
DFF_save_fm DFF_W5461(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31215));
DFF_save_fm DFF_W5462(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31225));
DFF_save_fm DFF_W5463(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31006));
DFF_save_fm DFF_W5464(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31016));
DFF_save_fm DFF_W5465(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31026));
DFF_save_fm DFF_W5466(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31106));
DFF_save_fm DFF_W5467(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31116));
DFF_save_fm DFF_W5468(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31126));
DFF_save_fm DFF_W5469(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31206));
DFF_save_fm DFF_W5470(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31216));
DFF_save_fm DFF_W5471(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31226));
DFF_save_fm DFF_W5472(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31007));
DFF_save_fm DFF_W5473(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31017));
DFF_save_fm DFF_W5474(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31027));
DFF_save_fm DFF_W5475(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31107));
DFF_save_fm DFF_W5476(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31117));
DFF_save_fm DFF_W5477(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31127));
DFF_save_fm DFF_W5478(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31207));
DFF_save_fm DFF_W5479(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31217));
DFF_save_fm DFF_W5480(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31227));
DFF_save_fm DFF_W5481(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31008));
DFF_save_fm DFF_W5482(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31018));
DFF_save_fm DFF_W5483(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31028));
DFF_save_fm DFF_W5484(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31108));
DFF_save_fm DFF_W5485(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31118));
DFF_save_fm DFF_W5486(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31128));
DFF_save_fm DFF_W5487(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31208));
DFF_save_fm DFF_W5488(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31218));
DFF_save_fm DFF_W5489(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31228));
DFF_save_fm DFF_W5490(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31009));
DFF_save_fm DFF_W5491(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31019));
DFF_save_fm DFF_W5492(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31029));
DFF_save_fm DFF_W5493(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31109));
DFF_save_fm DFF_W5494(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31119));
DFF_save_fm DFF_W5495(.clk(clk),.rstn(rstn),.reset_value(1),.q(W31129));
DFF_save_fm DFF_W5496(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31209));
DFF_save_fm DFF_W5497(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31219));
DFF_save_fm DFF_W5498(.clk(clk),.rstn(rstn),.reset_value(0),.q(W31229));
DFF_save_fm DFF_W5499(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3100A));
DFF_save_fm DFF_W5500(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3101A));
DFF_save_fm DFF_W5501(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3102A));
DFF_save_fm DFF_W5502(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3110A));
DFF_save_fm DFF_W5503(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3111A));
DFF_save_fm DFF_W5504(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3112A));
DFF_save_fm DFF_W5505(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120A));
DFF_save_fm DFF_W5506(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3121A));
DFF_save_fm DFF_W5507(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3122A));
DFF_save_fm DFF_W5508(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3100B));
DFF_save_fm DFF_W5509(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3101B));
DFF_save_fm DFF_W5510(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3102B));
DFF_save_fm DFF_W5511(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3110B));
DFF_save_fm DFF_W5512(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3111B));
DFF_save_fm DFF_W5513(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3112B));
DFF_save_fm DFF_W5514(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120B));
DFF_save_fm DFF_W5515(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3121B));
DFF_save_fm DFF_W5516(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3122B));
DFF_save_fm DFF_W5517(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3100C));
DFF_save_fm DFF_W5518(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3101C));
DFF_save_fm DFF_W5519(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3102C));
DFF_save_fm DFF_W5520(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3110C));
DFF_save_fm DFF_W5521(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3111C));
DFF_save_fm DFF_W5522(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3112C));
DFF_save_fm DFF_W5523(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120C));
DFF_save_fm DFF_W5524(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3121C));
DFF_save_fm DFF_W5525(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3122C));
DFF_save_fm DFF_W5526(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3100D));
DFF_save_fm DFF_W5527(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3101D));
DFF_save_fm DFF_W5528(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3102D));
DFF_save_fm DFF_W5529(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3110D));
DFF_save_fm DFF_W5530(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3111D));
DFF_save_fm DFF_W5531(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3112D));
DFF_save_fm DFF_W5532(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3120D));
DFF_save_fm DFF_W5533(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3121D));
DFF_save_fm DFF_W5534(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3122D));
DFF_save_fm DFF_W5535(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3100E));
DFF_save_fm DFF_W5536(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3101E));
DFF_save_fm DFF_W5537(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3102E));
DFF_save_fm DFF_W5538(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3110E));
DFF_save_fm DFF_W5539(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3111E));
DFF_save_fm DFF_W5540(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3112E));
DFF_save_fm DFF_W5541(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3120E));
DFF_save_fm DFF_W5542(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3121E));
DFF_save_fm DFF_W5543(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3122E));
DFF_save_fm DFF_W5544(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3100F));
DFF_save_fm DFF_W5545(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3101F));
DFF_save_fm DFF_W5546(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3102F));
DFF_save_fm DFF_W5547(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3110F));
DFF_save_fm DFF_W5548(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3111F));
DFF_save_fm DFF_W5549(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3112F));
DFF_save_fm DFF_W5550(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3120F));
DFF_save_fm DFF_W5551(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3121F));
DFF_save_fm DFF_W5552(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3122F));
DFF_save_fm DFF_W5553(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3100G));
DFF_save_fm DFF_W5554(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3101G));
DFF_save_fm DFF_W5555(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3102G));
DFF_save_fm DFF_W5556(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3110G));
DFF_save_fm DFF_W5557(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3111G));
DFF_save_fm DFF_W5558(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3112G));
DFF_save_fm DFF_W5559(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3120G));
DFF_save_fm DFF_W5560(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3121G));
DFF_save_fm DFF_W5561(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3122G));
DFF_save_fm DFF_W5562(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3100H));
DFF_save_fm DFF_W5563(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3101H));
DFF_save_fm DFF_W5564(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3102H));
DFF_save_fm DFF_W5565(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3110H));
DFF_save_fm DFF_W5566(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3111H));
DFF_save_fm DFF_W5567(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3112H));
DFF_save_fm DFF_W5568(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3120H));
DFF_save_fm DFF_W5569(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3121H));
DFF_save_fm DFF_W5570(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3122H));
DFF_save_fm DFF_W5571(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3100I));
DFF_save_fm DFF_W5572(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3101I));
DFF_save_fm DFF_W5573(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3102I));
DFF_save_fm DFF_W5574(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3110I));
DFF_save_fm DFF_W5575(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3111I));
DFF_save_fm DFF_W5576(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3112I));
DFF_save_fm DFF_W5577(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3120I));
DFF_save_fm DFF_W5578(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3121I));
DFF_save_fm DFF_W5579(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3122I));
DFF_save_fm DFF_W5580(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3100J));
DFF_save_fm DFF_W5581(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3101J));
DFF_save_fm DFF_W5582(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3102J));
DFF_save_fm DFF_W5583(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3110J));
DFF_save_fm DFF_W5584(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3111J));
DFF_save_fm DFF_W5585(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3112J));
DFF_save_fm DFF_W5586(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120J));
DFF_save_fm DFF_W5587(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3121J));
DFF_save_fm DFF_W5588(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3122J));
DFF_save_fm DFF_W5589(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3100K));
DFF_save_fm DFF_W5590(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3101K));
DFF_save_fm DFF_W5591(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3102K));
DFF_save_fm DFF_W5592(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3110K));
DFF_save_fm DFF_W5593(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3111K));
DFF_save_fm DFF_W5594(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3112K));
DFF_save_fm DFF_W5595(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120K));
DFF_save_fm DFF_W5596(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3121K));
DFF_save_fm DFF_W5597(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3122K));
DFF_save_fm DFF_W5598(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3100L));
DFF_save_fm DFF_W5599(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3101L));
DFF_save_fm DFF_W5600(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3102L));
DFF_save_fm DFF_W5601(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3110L));
DFF_save_fm DFF_W5602(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3111L));
DFF_save_fm DFF_W5603(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3112L));
DFF_save_fm DFF_W5604(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120L));
DFF_save_fm DFF_W5605(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3121L));
DFF_save_fm DFF_W5606(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3122L));
DFF_save_fm DFF_W5607(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3100M));
DFF_save_fm DFF_W5608(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3101M));
DFF_save_fm DFF_W5609(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3102M));
DFF_save_fm DFF_W5610(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3110M));
DFF_save_fm DFF_W5611(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3111M));
DFF_save_fm DFF_W5612(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3112M));
DFF_save_fm DFF_W5613(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120M));
DFF_save_fm DFF_W5614(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3121M));
DFF_save_fm DFF_W5615(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3122M));
DFF_save_fm DFF_W5616(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3100N));
DFF_save_fm DFF_W5617(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3101N));
DFF_save_fm DFF_W5618(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3102N));
DFF_save_fm DFF_W5619(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3110N));
DFF_save_fm DFF_W5620(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3111N));
DFF_save_fm DFF_W5621(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3112N));
DFF_save_fm DFF_W5622(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120N));
DFF_save_fm DFF_W5623(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3121N));
DFF_save_fm DFF_W5624(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3122N));
DFF_save_fm DFF_W5625(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3100O));
DFF_save_fm DFF_W5626(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3101O));
DFF_save_fm DFF_W5627(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3102O));
DFF_save_fm DFF_W5628(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3110O));
DFF_save_fm DFF_W5629(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3111O));
DFF_save_fm DFF_W5630(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3112O));
DFF_save_fm DFF_W5631(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120O));
DFF_save_fm DFF_W5632(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3121O));
DFF_save_fm DFF_W5633(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3122O));
DFF_save_fm DFF_W5634(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3100P));
DFF_save_fm DFF_W5635(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3101P));
DFF_save_fm DFF_W5636(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3102P));
DFF_save_fm DFF_W5637(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3110P));
DFF_save_fm DFF_W5638(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3111P));
DFF_save_fm DFF_W5639(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3112P));
DFF_save_fm DFF_W5640(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120P));
DFF_save_fm DFF_W5641(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3121P));
DFF_save_fm DFF_W5642(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3122P));
DFF_save_fm DFF_W5643(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3100Q));
DFF_save_fm DFF_W5644(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3101Q));
DFF_save_fm DFF_W5645(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3102Q));
DFF_save_fm DFF_W5646(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3110Q));
DFF_save_fm DFF_W5647(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3111Q));
DFF_save_fm DFF_W5648(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3112Q));
DFF_save_fm DFF_W5649(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120Q));
DFF_save_fm DFF_W5650(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3121Q));
DFF_save_fm DFF_W5651(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3122Q));
DFF_save_fm DFF_W5652(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3100R));
DFF_save_fm DFF_W5653(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3101R));
DFF_save_fm DFF_W5654(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3102R));
DFF_save_fm DFF_W5655(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3110R));
DFF_save_fm DFF_W5656(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3111R));
DFF_save_fm DFF_W5657(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3112R));
DFF_save_fm DFF_W5658(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120R));
DFF_save_fm DFF_W5659(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3121R));
DFF_save_fm DFF_W5660(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3122R));
DFF_save_fm DFF_W5661(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3100S));
DFF_save_fm DFF_W5662(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3101S));
DFF_save_fm DFF_W5663(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3102S));
DFF_save_fm DFF_W5664(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3110S));
DFF_save_fm DFF_W5665(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3111S));
DFF_save_fm DFF_W5666(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3112S));
DFF_save_fm DFF_W5667(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120S));
DFF_save_fm DFF_W5668(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3121S));
DFF_save_fm DFF_W5669(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3122S));
DFF_save_fm DFF_W5670(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3100T));
DFF_save_fm DFF_W5671(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3101T));
DFF_save_fm DFF_W5672(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3102T));
DFF_save_fm DFF_W5673(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3110T));
DFF_save_fm DFF_W5674(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3111T));
DFF_save_fm DFF_W5675(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3112T));
DFF_save_fm DFF_W5676(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120T));
DFF_save_fm DFF_W5677(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3121T));
DFF_save_fm DFF_W5678(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3122T));
DFF_save_fm DFF_W5679(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3100U));
DFF_save_fm DFF_W5680(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3101U));
DFF_save_fm DFF_W5681(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3102U));
DFF_save_fm DFF_W5682(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3110U));
DFF_save_fm DFF_W5683(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3111U));
DFF_save_fm DFF_W5684(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3112U));
DFF_save_fm DFF_W5685(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120U));
DFF_save_fm DFF_W5686(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3121U));
DFF_save_fm DFF_W5687(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3122U));
DFF_save_fm DFF_W5688(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3100V));
DFF_save_fm DFF_W5689(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3101V));
DFF_save_fm DFF_W5690(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3102V));
DFF_save_fm DFF_W5691(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3110V));
DFF_save_fm DFF_W5692(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3111V));
DFF_save_fm DFF_W5693(.clk(clk),.rstn(rstn),.reset_value(0),.q(W3112V));
DFF_save_fm DFF_W5694(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3120V));
DFF_save_fm DFF_W5695(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3121V));
DFF_save_fm DFF_W5696(.clk(clk),.rstn(rstn),.reset_value(1),.q(W3122V));
ninexnine_unit ninexnine_unit_7572(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W30000),
				.b1(W30010),
				.b2(W30020),
				.b3(W30100),
				.b4(W30110),
				.b5(W30120),
				.b6(W30200),
				.b7(W30210),
				.b8(W30220),
				.c(c30000)
);

ninexnine_unit ninexnine_unit_7573(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W30001),
				.b1(W30011),
				.b2(W30021),
				.b3(W30101),
				.b4(W30111),
				.b5(W30121),
				.b6(W30201),
				.b7(W30211),
				.b8(W30221),
				.c(c31000)
);

ninexnine_unit ninexnine_unit_7574(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W30002),
				.b1(W30012),
				.b2(W30022),
				.b3(W30102),
				.b4(W30112),
				.b5(W30122),
				.b6(W30202),
				.b7(W30212),
				.b8(W30222),
				.c(c32000)
);

ninexnine_unit ninexnine_unit_7575(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W30003),
				.b1(W30013),
				.b2(W30023),
				.b3(W30103),
				.b4(W30113),
				.b5(W30123),
				.b6(W30203),
				.b7(W30213),
				.b8(W30223),
				.c(c33000)
);

ninexnine_unit ninexnine_unit_7576(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W30004),
				.b1(W30014),
				.b2(W30024),
				.b3(W30104),
				.b4(W30114),
				.b5(W30124),
				.b6(W30204),
				.b7(W30214),
				.b8(W30224),
				.c(c34000)
);

ninexnine_unit ninexnine_unit_7577(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W30005),
				.b1(W30015),
				.b2(W30025),
				.b3(W30105),
				.b4(W30115),
				.b5(W30125),
				.b6(W30205),
				.b7(W30215),
				.b8(W30225),
				.c(c35000)
);

ninexnine_unit ninexnine_unit_7578(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W30006),
				.b1(W30016),
				.b2(W30026),
				.b3(W30106),
				.b4(W30116),
				.b5(W30126),
				.b6(W30206),
				.b7(W30216),
				.b8(W30226),
				.c(c36000)
);

ninexnine_unit ninexnine_unit_7579(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W30007),
				.b1(W30017),
				.b2(W30027),
				.b3(W30107),
				.b4(W30117),
				.b5(W30127),
				.b6(W30207),
				.b7(W30217),
				.b8(W30227),
				.c(c37000)
);

ninexnine_unit ninexnine_unit_7580(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W30008),
				.b1(W30018),
				.b2(W30028),
				.b3(W30108),
				.b4(W30118),
				.b5(W30128),
				.b6(W30208),
				.b7(W30218),
				.b8(W30228),
				.c(c38000)
);

ninexnine_unit ninexnine_unit_7581(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W30009),
				.b1(W30019),
				.b2(W30029),
				.b3(W30109),
				.b4(W30119),
				.b5(W30129),
				.b6(W30209),
				.b7(W30219),
				.b8(W30229),
				.c(c39000)
);

ninexnine_unit ninexnine_unit_7582(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3000A),
				.b1(W3001A),
				.b2(W3002A),
				.b3(W3010A),
				.b4(W3011A),
				.b5(W3012A),
				.b6(W3020A),
				.b7(W3021A),
				.b8(W3022A),
				.c(c3A000)
);

ninexnine_unit ninexnine_unit_7583(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3000B),
				.b1(W3001B),
				.b2(W3002B),
				.b3(W3010B),
				.b4(W3011B),
				.b5(W3012B),
				.b6(W3020B),
				.b7(W3021B),
				.b8(W3022B),
				.c(c3B000)
);

ninexnine_unit ninexnine_unit_7584(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3000C),
				.b1(W3001C),
				.b2(W3002C),
				.b3(W3010C),
				.b4(W3011C),
				.b5(W3012C),
				.b6(W3020C),
				.b7(W3021C),
				.b8(W3022C),
				.c(c3C000)
);

ninexnine_unit ninexnine_unit_7585(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3000D),
				.b1(W3001D),
				.b2(W3002D),
				.b3(W3010D),
				.b4(W3011D),
				.b5(W3012D),
				.b6(W3020D),
				.b7(W3021D),
				.b8(W3022D),
				.c(c3D000)
);

ninexnine_unit ninexnine_unit_7586(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3000E),
				.b1(W3001E),
				.b2(W3002E),
				.b3(W3010E),
				.b4(W3011E),
				.b5(W3012E),
				.b6(W3020E),
				.b7(W3021E),
				.b8(W3022E),
				.c(c3E000)
);

ninexnine_unit ninexnine_unit_7587(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3000F),
				.b1(W3001F),
				.b2(W3002F),
				.b3(W3010F),
				.b4(W3011F),
				.b5(W3012F),
				.b6(W3020F),
				.b7(W3021F),
				.b8(W3022F),
				.c(c3F000)
);

ninexnine_unit ninexnine_unit_7588(
				.clk(clk),
				.rstn(rstn),
				.a0(P300G),
				.a1(P301G),
				.a2(P302G),
				.a3(P310G),
				.a4(P311G),
				.a5(P312G),
				.a6(P320G),
				.a7(P321G),
				.a8(P322G),
				.b0(W3000G),
				.b1(W3001G),
				.b2(W3002G),
				.b3(W3010G),
				.b4(W3011G),
				.b5(W3012G),
				.b6(W3020G),
				.b7(W3021G),
				.b8(W3022G),
				.c(c3G000)
);

ninexnine_unit ninexnine_unit_7589(
				.clk(clk),
				.rstn(rstn),
				.a0(P300H),
				.a1(P301H),
				.a2(P302H),
				.a3(P310H),
				.a4(P311H),
				.a5(P312H),
				.a6(P320H),
				.a7(P321H),
				.a8(P322H),
				.b0(W3000H),
				.b1(W3001H),
				.b2(W3002H),
				.b3(W3010H),
				.b4(W3011H),
				.b5(W3012H),
				.b6(W3020H),
				.b7(W3021H),
				.b8(W3022H),
				.c(c3H000)
);

ninexnine_unit ninexnine_unit_7590(
				.clk(clk),
				.rstn(rstn),
				.a0(P300I),
				.a1(P301I),
				.a2(P302I),
				.a3(P310I),
				.a4(P311I),
				.a5(P312I),
				.a6(P320I),
				.a7(P321I),
				.a8(P322I),
				.b0(W3000I),
				.b1(W3001I),
				.b2(W3002I),
				.b3(W3010I),
				.b4(W3011I),
				.b5(W3012I),
				.b6(W3020I),
				.b7(W3021I),
				.b8(W3022I),
				.c(c3I000)
);

ninexnine_unit ninexnine_unit_7591(
				.clk(clk),
				.rstn(rstn),
				.a0(P300J),
				.a1(P301J),
				.a2(P302J),
				.a3(P310J),
				.a4(P311J),
				.a5(P312J),
				.a6(P320J),
				.a7(P321J),
				.a8(P322J),
				.b0(W3000J),
				.b1(W3001J),
				.b2(W3002J),
				.b3(W3010J),
				.b4(W3011J),
				.b5(W3012J),
				.b6(W3020J),
				.b7(W3021J),
				.b8(W3022J),
				.c(c3J000)
);

ninexnine_unit ninexnine_unit_7592(
				.clk(clk),
				.rstn(rstn),
				.a0(P300K),
				.a1(P301K),
				.a2(P302K),
				.a3(P310K),
				.a4(P311K),
				.a5(P312K),
				.a6(P320K),
				.a7(P321K),
				.a8(P322K),
				.b0(W3000K),
				.b1(W3001K),
				.b2(W3002K),
				.b3(W3010K),
				.b4(W3011K),
				.b5(W3012K),
				.b6(W3020K),
				.b7(W3021K),
				.b8(W3022K),
				.c(c3K000)
);

ninexnine_unit ninexnine_unit_7593(
				.clk(clk),
				.rstn(rstn),
				.a0(P300L),
				.a1(P301L),
				.a2(P302L),
				.a3(P310L),
				.a4(P311L),
				.a5(P312L),
				.a6(P320L),
				.a7(P321L),
				.a8(P322L),
				.b0(W3000L),
				.b1(W3001L),
				.b2(W3002L),
				.b3(W3010L),
				.b4(W3011L),
				.b5(W3012L),
				.b6(W3020L),
				.b7(W3021L),
				.b8(W3022L),
				.c(c3L000)
);

ninexnine_unit ninexnine_unit_7594(
				.clk(clk),
				.rstn(rstn),
				.a0(P300M),
				.a1(P301M),
				.a2(P302M),
				.a3(P310M),
				.a4(P311M),
				.a5(P312M),
				.a6(P320M),
				.a7(P321M),
				.a8(P322M),
				.b0(W3000M),
				.b1(W3001M),
				.b2(W3002M),
				.b3(W3010M),
				.b4(W3011M),
				.b5(W3012M),
				.b6(W3020M),
				.b7(W3021M),
				.b8(W3022M),
				.c(c3M000)
);

ninexnine_unit ninexnine_unit_7595(
				.clk(clk),
				.rstn(rstn),
				.a0(P300N),
				.a1(P301N),
				.a2(P302N),
				.a3(P310N),
				.a4(P311N),
				.a5(P312N),
				.a6(P320N),
				.a7(P321N),
				.a8(P322N),
				.b0(W3000N),
				.b1(W3001N),
				.b2(W3002N),
				.b3(W3010N),
				.b4(W3011N),
				.b5(W3012N),
				.b6(W3020N),
				.b7(W3021N),
				.b8(W3022N),
				.c(c3N000)
);

ninexnine_unit ninexnine_unit_7596(
				.clk(clk),
				.rstn(rstn),
				.a0(P300O),
				.a1(P301O),
				.a2(P302O),
				.a3(P310O),
				.a4(P311O),
				.a5(P312O),
				.a6(P320O),
				.a7(P321O),
				.a8(P322O),
				.b0(W3000O),
				.b1(W3001O),
				.b2(W3002O),
				.b3(W3010O),
				.b4(W3011O),
				.b5(W3012O),
				.b6(W3020O),
				.b7(W3021O),
				.b8(W3022O),
				.c(c3O000)
);

ninexnine_unit ninexnine_unit_7597(
				.clk(clk),
				.rstn(rstn),
				.a0(P300P),
				.a1(P301P),
				.a2(P302P),
				.a3(P310P),
				.a4(P311P),
				.a5(P312P),
				.a6(P320P),
				.a7(P321P),
				.a8(P322P),
				.b0(W3000P),
				.b1(W3001P),
				.b2(W3002P),
				.b3(W3010P),
				.b4(W3011P),
				.b5(W3012P),
				.b6(W3020P),
				.b7(W3021P),
				.b8(W3022P),
				.c(c3P000)
);

ninexnine_unit ninexnine_unit_7598(
				.clk(clk),
				.rstn(rstn),
				.a0(P300Q),
				.a1(P301Q),
				.a2(P302Q),
				.a3(P310Q),
				.a4(P311Q),
				.a5(P312Q),
				.a6(P320Q),
				.a7(P321Q),
				.a8(P322Q),
				.b0(W3000Q),
				.b1(W3001Q),
				.b2(W3002Q),
				.b3(W3010Q),
				.b4(W3011Q),
				.b5(W3012Q),
				.b6(W3020Q),
				.b7(W3021Q),
				.b8(W3022Q),
				.c(c3Q000)
);

ninexnine_unit ninexnine_unit_7599(
				.clk(clk),
				.rstn(rstn),
				.a0(P300R),
				.a1(P301R),
				.a2(P302R),
				.a3(P310R),
				.a4(P311R),
				.a5(P312R),
				.a6(P320R),
				.a7(P321R),
				.a8(P322R),
				.b0(W3000R),
				.b1(W3001R),
				.b2(W3002R),
				.b3(W3010R),
				.b4(W3011R),
				.b5(W3012R),
				.b6(W3020R),
				.b7(W3021R),
				.b8(W3022R),
				.c(c3R000)
);

ninexnine_unit ninexnine_unit_7600(
				.clk(clk),
				.rstn(rstn),
				.a0(P300S),
				.a1(P301S),
				.a2(P302S),
				.a3(P310S),
				.a4(P311S),
				.a5(P312S),
				.a6(P320S),
				.a7(P321S),
				.a8(P322S),
				.b0(W3000S),
				.b1(W3001S),
				.b2(W3002S),
				.b3(W3010S),
				.b4(W3011S),
				.b5(W3012S),
				.b6(W3020S),
				.b7(W3021S),
				.b8(W3022S),
				.c(c3S000)
);

ninexnine_unit ninexnine_unit_7601(
				.clk(clk),
				.rstn(rstn),
				.a0(P300T),
				.a1(P301T),
				.a2(P302T),
				.a3(P310T),
				.a4(P311T),
				.a5(P312T),
				.a6(P320T),
				.a7(P321T),
				.a8(P322T),
				.b0(W3000T),
				.b1(W3001T),
				.b2(W3002T),
				.b3(W3010T),
				.b4(W3011T),
				.b5(W3012T),
				.b6(W3020T),
				.b7(W3021T),
				.b8(W3022T),
				.c(c3T000)
);

ninexnine_unit ninexnine_unit_7602(
				.clk(clk),
				.rstn(rstn),
				.a0(P300U),
				.a1(P301U),
				.a2(P302U),
				.a3(P310U),
				.a4(P311U),
				.a5(P312U),
				.a6(P320U),
				.a7(P321U),
				.a8(P322U),
				.b0(W3000U),
				.b1(W3001U),
				.b2(W3002U),
				.b3(W3010U),
				.b4(W3011U),
				.b5(W3012U),
				.b6(W3020U),
				.b7(W3021U),
				.b8(W3022U),
				.c(c3U000)
);

ninexnine_unit ninexnine_unit_7603(
				.clk(clk),
				.rstn(rstn),
				.a0(P300V),
				.a1(P301V),
				.a2(P302V),
				.a3(P310V),
				.a4(P311V),
				.a5(P312V),
				.a6(P320V),
				.a7(P321V),
				.a8(P322V),
				.b0(W3000V),
				.b1(W3001V),
				.b2(W3002V),
				.b3(W3010V),
				.b4(W3011V),
				.b5(W3012V),
				.b6(W3020V),
				.b7(W3021V),
				.b8(W3022V),
				.c(c3V000)
);

assign C3000=c30000+c31000+c32000+c33000+c34000+c35000+c36000+c37000+c38000+c39000+c3A000+c3B000+c3C000+c3D000+c3E000+c3F000+c3G000+c3H000+c3I000+c3J000+c3K000+c3L000+c3M000+c3N000+c3O000+c3P000+c3Q000+c3R000+c3S000+c3T000+c3U000+c3V000;
assign A3000=(C3000>=0)?1:0;

assign P4000=A3000;

ninexnine_unit ninexnine_unit_7604(
				.clk(clk),
				.rstn(rstn),
				.a0(P3000),
				.a1(P3010),
				.a2(P3020),
				.a3(P3100),
				.a4(P3110),
				.a5(P3120),
				.a6(P3200),
				.a7(P3210),
				.a8(P3220),
				.b0(W31000),
				.b1(W31010),
				.b2(W31020),
				.b3(W31100),
				.b4(W31110),
				.b5(W31120),
				.b6(W31200),
				.b7(W31210),
				.b8(W31220),
				.c(c30001)
);

ninexnine_unit ninexnine_unit_7605(
				.clk(clk),
				.rstn(rstn),
				.a0(P3001),
				.a1(P3011),
				.a2(P3021),
				.a3(P3101),
				.a4(P3111),
				.a5(P3121),
				.a6(P3201),
				.a7(P3211),
				.a8(P3221),
				.b0(W31001),
				.b1(W31011),
				.b2(W31021),
				.b3(W31101),
				.b4(W31111),
				.b5(W31121),
				.b6(W31201),
				.b7(W31211),
				.b8(W31221),
				.c(c31001)
);

ninexnine_unit ninexnine_unit_7606(
				.clk(clk),
				.rstn(rstn),
				.a0(P3002),
				.a1(P3012),
				.a2(P3022),
				.a3(P3102),
				.a4(P3112),
				.a5(P3122),
				.a6(P3202),
				.a7(P3212),
				.a8(P3222),
				.b0(W31002),
				.b1(W31012),
				.b2(W31022),
				.b3(W31102),
				.b4(W31112),
				.b5(W31122),
				.b6(W31202),
				.b7(W31212),
				.b8(W31222),
				.c(c32001)
);

ninexnine_unit ninexnine_unit_7607(
				.clk(clk),
				.rstn(rstn),
				.a0(P3003),
				.a1(P3013),
				.a2(P3023),
				.a3(P3103),
				.a4(P3113),
				.a5(P3123),
				.a6(P3203),
				.a7(P3213),
				.a8(P3223),
				.b0(W31003),
				.b1(W31013),
				.b2(W31023),
				.b3(W31103),
				.b4(W31113),
				.b5(W31123),
				.b6(W31203),
				.b7(W31213),
				.b8(W31223),
				.c(c33001)
);

ninexnine_unit ninexnine_unit_7608(
				.clk(clk),
				.rstn(rstn),
				.a0(P3004),
				.a1(P3014),
				.a2(P3024),
				.a3(P3104),
				.a4(P3114),
				.a5(P3124),
				.a6(P3204),
				.a7(P3214),
				.a8(P3224),
				.b0(W31004),
				.b1(W31014),
				.b2(W31024),
				.b3(W31104),
				.b4(W31114),
				.b5(W31124),
				.b6(W31204),
				.b7(W31214),
				.b8(W31224),
				.c(c34001)
);

ninexnine_unit ninexnine_unit_7609(
				.clk(clk),
				.rstn(rstn),
				.a0(P3005),
				.a1(P3015),
				.a2(P3025),
				.a3(P3105),
				.a4(P3115),
				.a5(P3125),
				.a6(P3205),
				.a7(P3215),
				.a8(P3225),
				.b0(W31005),
				.b1(W31015),
				.b2(W31025),
				.b3(W31105),
				.b4(W31115),
				.b5(W31125),
				.b6(W31205),
				.b7(W31215),
				.b8(W31225),
				.c(c35001)
);

ninexnine_unit ninexnine_unit_7610(
				.clk(clk),
				.rstn(rstn),
				.a0(P3006),
				.a1(P3016),
				.a2(P3026),
				.a3(P3106),
				.a4(P3116),
				.a5(P3126),
				.a6(P3206),
				.a7(P3216),
				.a8(P3226),
				.b0(W31006),
				.b1(W31016),
				.b2(W31026),
				.b3(W31106),
				.b4(W31116),
				.b5(W31126),
				.b6(W31206),
				.b7(W31216),
				.b8(W31226),
				.c(c36001)
);

ninexnine_unit ninexnine_unit_7611(
				.clk(clk),
				.rstn(rstn),
				.a0(P3007),
				.a1(P3017),
				.a2(P3027),
				.a3(P3107),
				.a4(P3117),
				.a5(P3127),
				.a6(P3207),
				.a7(P3217),
				.a8(P3227),
				.b0(W31007),
				.b1(W31017),
				.b2(W31027),
				.b3(W31107),
				.b4(W31117),
				.b5(W31127),
				.b6(W31207),
				.b7(W31217),
				.b8(W31227),
				.c(c37001)
);

ninexnine_unit ninexnine_unit_7612(
				.clk(clk),
				.rstn(rstn),
				.a0(P3008),
				.a1(P3018),
				.a2(P3028),
				.a3(P3108),
				.a4(P3118),
				.a5(P3128),
				.a6(P3208),
				.a7(P3218),
				.a8(P3228),
				.b0(W31008),
				.b1(W31018),
				.b2(W31028),
				.b3(W31108),
				.b4(W31118),
				.b5(W31128),
				.b6(W31208),
				.b7(W31218),
				.b8(W31228),
				.c(c38001)
);

ninexnine_unit ninexnine_unit_7613(
				.clk(clk),
				.rstn(rstn),
				.a0(P3009),
				.a1(P3019),
				.a2(P3029),
				.a3(P3109),
				.a4(P3119),
				.a5(P3129),
				.a6(P3209),
				.a7(P3219),
				.a8(P3229),
				.b0(W31009),
				.b1(W31019),
				.b2(W31029),
				.b3(W31109),
				.b4(W31119),
				.b5(W31129),
				.b6(W31209),
				.b7(W31219),
				.b8(W31229),
				.c(c39001)
);

ninexnine_unit ninexnine_unit_7614(
				.clk(clk),
				.rstn(rstn),
				.a0(P300A),
				.a1(P301A),
				.a2(P302A),
				.a3(P310A),
				.a4(P311A),
				.a5(P312A),
				.a6(P320A),
				.a7(P321A),
				.a8(P322A),
				.b0(W3100A),
				.b1(W3101A),
				.b2(W3102A),
				.b3(W3110A),
				.b4(W3111A),
				.b5(W3112A),
				.b6(W3120A),
				.b7(W3121A),
				.b8(W3122A),
				.c(c3A001)
);

ninexnine_unit ninexnine_unit_7615(
				.clk(clk),
				.rstn(rstn),
				.a0(P300B),
				.a1(P301B),
				.a2(P302B),
				.a3(P310B),
				.a4(P311B),
				.a5(P312B),
				.a6(P320B),
				.a7(P321B),
				.a8(P322B),
				.b0(W3100B),
				.b1(W3101B),
				.b2(W3102B),
				.b3(W3110B),
				.b4(W3111B),
				.b5(W3112B),
				.b6(W3120B),
				.b7(W3121B),
				.b8(W3122B),
				.c(c3B001)
);

ninexnine_unit ninexnine_unit_7616(
				.clk(clk),
				.rstn(rstn),
				.a0(P300C),
				.a1(P301C),
				.a2(P302C),
				.a3(P310C),
				.a4(P311C),
				.a5(P312C),
				.a6(P320C),
				.a7(P321C),
				.a8(P322C),
				.b0(W3100C),
				.b1(W3101C),
				.b2(W3102C),
				.b3(W3110C),
				.b4(W3111C),
				.b5(W3112C),
				.b6(W3120C),
				.b7(W3121C),
				.b8(W3122C),
				.c(c3C001)
);

ninexnine_unit ninexnine_unit_7617(
				.clk(clk),
				.rstn(rstn),
				.a0(P300D),
				.a1(P301D),
				.a2(P302D),
				.a3(P310D),
				.a4(P311D),
				.a5(P312D),
				.a6(P320D),
				.a7(P321D),
				.a8(P322D),
				.b0(W3100D),
				.b1(W3101D),
				.b2(W3102D),
				.b3(W3110D),
				.b4(W3111D),
				.b5(W3112D),
				.b6(W3120D),
				.b7(W3121D),
				.b8(W3122D),
				.c(c3D001)
);

ninexnine_unit ninexnine_unit_7618(
				.clk(clk),
				.rstn(rstn),
				.a0(P300E),
				.a1(P301E),
				.a2(P302E),
				.a3(P310E),
				.a4(P311E),
				.a5(P312E),
				.a6(P320E),
				.a7(P321E),
				.a8(P322E),
				.b0(W3100E),
				.b1(W3101E),
				.b2(W3102E),
				.b3(W3110E),
				.b4(W3111E),
				.b5(W3112E),
				.b6(W3120E),
				.b7(W3121E),
				.b8(W3122E),
				.c(c3E001)
);

ninexnine_unit ninexnine_unit_7619(
				.clk(clk),
				.rstn(rstn),
				.a0(P300F),
				.a1(P301F),
				.a2(P302F),
				.a3(P310F),
				.a4(P311F),
				.a5(P312F),
				.a6(P320F),
				.a7(P321F),
				.a8(P322F),
				.b0(W3100F),
				.b1(W3101F),
				.b2(W3102F),
				.b3(W3110F),
				.b4(W3111F),
				.b5(W3112F),
				.b6(W3120F),
				.b7(W3121F),
				.b8(W3122F),
				.c(c3F001)
);

ninexnine_unit ninexnine_unit_7620(
				.clk(clk),
				.rstn(rstn),
				.a0(P300G),
				.a1(P301G),
				.a2(P302G),
				.a3(P310G),
				.a4(P311G),
				.a5(P312G),
				.a6(P320G),
				.a7(P321G),
				.a8(P322G),
				.b0(W3100G),
				.b1(W3101G),
				.b2(W3102G),
				.b3(W3110G),
				.b4(W3111G),
				.b5(W3112G),
				.b6(W3120G),
				.b7(W3121G),
				.b8(W3122G),
				.c(c3G001)
);

ninexnine_unit ninexnine_unit_7621(
				.clk(clk),
				.rstn(rstn),
				.a0(P300H),
				.a1(P301H),
				.a2(P302H),
				.a3(P310H),
				.a4(P311H),
				.a5(P312H),
				.a6(P320H),
				.a7(P321H),
				.a8(P322H),
				.b0(W3100H),
				.b1(W3101H),
				.b2(W3102H),
				.b3(W3110H),
				.b4(W3111H),
				.b5(W3112H),
				.b6(W3120H),
				.b7(W3121H),
				.b8(W3122H),
				.c(c3H001)
);

ninexnine_unit ninexnine_unit_7622(
				.clk(clk),
				.rstn(rstn),
				.a0(P300I),
				.a1(P301I),
				.a2(P302I),
				.a3(P310I),
				.a4(P311I),
				.a5(P312I),
				.a6(P320I),
				.a7(P321I),
				.a8(P322I),
				.b0(W3100I),
				.b1(W3101I),
				.b2(W3102I),
				.b3(W3110I),
				.b4(W3111I),
				.b5(W3112I),
				.b6(W3120I),
				.b7(W3121I),
				.b8(W3122I),
				.c(c3I001)
);

ninexnine_unit ninexnine_unit_7623(
				.clk(clk),
				.rstn(rstn),
				.a0(P300J),
				.a1(P301J),
				.a2(P302J),
				.a3(P310J),
				.a4(P311J),
				.a5(P312J),
				.a6(P320J),
				.a7(P321J),
				.a8(P322J),
				.b0(W3100J),
				.b1(W3101J),
				.b2(W3102J),
				.b3(W3110J),
				.b4(W3111J),
				.b5(W3112J),
				.b6(W3120J),
				.b7(W3121J),
				.b8(W3122J),
				.c(c3J001)
);

ninexnine_unit ninexnine_unit_7624(
				.clk(clk),
				.rstn(rstn),
				.a0(P300K),
				.a1(P301K),
				.a2(P302K),
				.a3(P310K),
				.a4(P311K),
				.a5(P312K),
				.a6(P320K),
				.a7(P321K),
				.a8(P322K),
				.b0(W3100K),
				.b1(W3101K),
				.b2(W3102K),
				.b3(W3110K),
				.b4(W3111K),
				.b5(W3112K),
				.b6(W3120K),
				.b7(W3121K),
				.b8(W3122K),
				.c(c3K001)
);

ninexnine_unit ninexnine_unit_7625(
				.clk(clk),
				.rstn(rstn),
				.a0(P300L),
				.a1(P301L),
				.a2(P302L),
				.a3(P310L),
				.a4(P311L),
				.a5(P312L),
				.a6(P320L),
				.a7(P321L),
				.a8(P322L),
				.b0(W3100L),
				.b1(W3101L),
				.b2(W3102L),
				.b3(W3110L),
				.b4(W3111L),
				.b5(W3112L),
				.b6(W3120L),
				.b7(W3121L),
				.b8(W3122L),
				.c(c3L001)
);

ninexnine_unit ninexnine_unit_7626(
				.clk(clk),
				.rstn(rstn),
				.a0(P300M),
				.a1(P301M),
				.a2(P302M),
				.a3(P310M),
				.a4(P311M),
				.a5(P312M),
				.a6(P320M),
				.a7(P321M),
				.a8(P322M),
				.b0(W3100M),
				.b1(W3101M),
				.b2(W3102M),
				.b3(W3110M),
				.b4(W3111M),
				.b5(W3112M),
				.b6(W3120M),
				.b7(W3121M),
				.b8(W3122M),
				.c(c3M001)
);

ninexnine_unit ninexnine_unit_7627(
				.clk(clk),
				.rstn(rstn),
				.a0(P300N),
				.a1(P301N),
				.a2(P302N),
				.a3(P310N),
				.a4(P311N),
				.a5(P312N),
				.a6(P320N),
				.a7(P321N),
				.a8(P322N),
				.b0(W3100N),
				.b1(W3101N),
				.b2(W3102N),
				.b3(W3110N),
				.b4(W3111N),
				.b5(W3112N),
				.b6(W3120N),
				.b7(W3121N),
				.b8(W3122N),
				.c(c3N001)
);

ninexnine_unit ninexnine_unit_7628(
				.clk(clk),
				.rstn(rstn),
				.a0(P300O),
				.a1(P301O),
				.a2(P302O),
				.a3(P310O),
				.a4(P311O),
				.a5(P312O),
				.a6(P320O),
				.a7(P321O),
				.a8(P322O),
				.b0(W3100O),
				.b1(W3101O),
				.b2(W3102O),
				.b3(W3110O),
				.b4(W3111O),
				.b5(W3112O),
				.b6(W3120O),
				.b7(W3121O),
				.b8(W3122O),
				.c(c3O001)
);

ninexnine_unit ninexnine_unit_7629(
				.clk(clk),
				.rstn(rstn),
				.a0(P300P),
				.a1(P301P),
				.a2(P302P),
				.a3(P310P),
				.a4(P311P),
				.a5(P312P),
				.a6(P320P),
				.a7(P321P),
				.a8(P322P),
				.b0(W3100P),
				.b1(W3101P),
				.b2(W3102P),
				.b3(W3110P),
				.b4(W3111P),
				.b5(W3112P),
				.b6(W3120P),
				.b7(W3121P),
				.b8(W3122P),
				.c(c3P001)
);

ninexnine_unit ninexnine_unit_7630(
				.clk(clk),
				.rstn(rstn),
				.a0(P300Q),
				.a1(P301Q),
				.a2(P302Q),
				.a3(P310Q),
				.a4(P311Q),
				.a5(P312Q),
				.a6(P320Q),
				.a7(P321Q),
				.a8(P322Q),
				.b0(W3100Q),
				.b1(W3101Q),
				.b2(W3102Q),
				.b3(W3110Q),
				.b4(W3111Q),
				.b5(W3112Q),
				.b6(W3120Q),
				.b7(W3121Q),
				.b8(W3122Q),
				.c(c3Q001)
);

ninexnine_unit ninexnine_unit_7631(
				.clk(clk),
				.rstn(rstn),
				.a0(P300R),
				.a1(P301R),
				.a2(P302R),
				.a3(P310R),
				.a4(P311R),
				.a5(P312R),
				.a6(P320R),
				.a7(P321R),
				.a8(P322R),
				.b0(W3100R),
				.b1(W3101R),
				.b2(W3102R),
				.b3(W3110R),
				.b4(W3111R),
				.b5(W3112R),
				.b6(W3120R),
				.b7(W3121R),
				.b8(W3122R),
				.c(c3R001)
);

ninexnine_unit ninexnine_unit_7632(
				.clk(clk),
				.rstn(rstn),
				.a0(P300S),
				.a1(P301S),
				.a2(P302S),
				.a3(P310S),
				.a4(P311S),
				.a5(P312S),
				.a6(P320S),
				.a7(P321S),
				.a8(P322S),
				.b0(W3100S),
				.b1(W3101S),
				.b2(W3102S),
				.b3(W3110S),
				.b4(W3111S),
				.b5(W3112S),
				.b6(W3120S),
				.b7(W3121S),
				.b8(W3122S),
				.c(c3S001)
);

ninexnine_unit ninexnine_unit_7633(
				.clk(clk),
				.rstn(rstn),
				.a0(P300T),
				.a1(P301T),
				.a2(P302T),
				.a3(P310T),
				.a4(P311T),
				.a5(P312T),
				.a6(P320T),
				.a7(P321T),
				.a8(P322T),
				.b0(W3100T),
				.b1(W3101T),
				.b2(W3102T),
				.b3(W3110T),
				.b4(W3111T),
				.b5(W3112T),
				.b6(W3120T),
				.b7(W3121T),
				.b8(W3122T),
				.c(c3T001)
);

ninexnine_unit ninexnine_unit_7634(
				.clk(clk),
				.rstn(rstn),
				.a0(P300U),
				.a1(P301U),
				.a2(P302U),
				.a3(P310U),
				.a4(P311U),
				.a5(P312U),
				.a6(P320U),
				.a7(P321U),
				.a8(P322U),
				.b0(W3100U),
				.b1(W3101U),
				.b2(W3102U),
				.b3(W3110U),
				.b4(W3111U),
				.b5(W3112U),
				.b6(W3120U),
				.b7(W3121U),
				.b8(W3122U),
				.c(c3U001)
);

ninexnine_unit ninexnine_unit_7635(
				.clk(clk),
				.rstn(rstn),
				.a0(P300V),
				.a1(P301V),
				.a2(P302V),
				.a3(P310V),
				.a4(P311V),
				.a5(P312V),
				.a6(P320V),
				.a7(P321V),
				.a8(P322V),
				.b0(W3100V),
				.b1(W3101V),
				.b2(W3102V),
				.b3(W3110V),
				.b4(W3111V),
				.b5(W3112V),
				.b6(W3120V),
				.b7(W3121V),
				.b8(W3122V),
				.c(c3V001)
);

assign C3001=c30001+c31001+c32001+c33001+c34001+c35001+c36001+c37001+c38001+c39001+c3A001+c3B001+c3C001+c3D001+c3E001+c3F001+c3G001+c3H001+c3I001+c3J001+c3K001+c3L001+c3M001+c3N001+c3O001+c3P001+c3Q001+c3R001+c3S001+c3T001+c3U001+c3V001;
assign A3001=(C3001>=0)?1:0;

assign P4001=A3001;

endmodule
//layer4 done, begain next layer
