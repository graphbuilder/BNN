module tb_test_layer0(

);
reg clk,rstn;
test_layer0 test_layer0(
clk,
rstn
);
reg mem[14*14*4-1:0];
always #5 clk=~clk;
initial
begin
clk=0;
rstn=0;
$readmemb("D:/work/PROJ_5/proj_2/src/to_csma/test_tb/answer_layer_0.txt",mem);
#10;
rstn=1;
end
reg [31:0]count;
always@(posedge clk or negedge rstn)
	if(~rstn)
		count<=0;
	else
		count<=count+1;

reg Pass_0;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_0<=0;
	else if(count>=2)
		begin
			if(tb_test_layer0.test_layer0.P1110==mem[0])
				Pass_0<=1;
			else
				Pass_0<=0;
		end

reg Pass_1;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_1<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1120==mem[1])&&(Pass_0))
				Pass_1<=1;
			else
				Pass_1<=0;
		end

reg Pass_2;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_2<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1130==mem[2])&&(Pass_1))
				Pass_2<=1;
			else
				Pass_2<=0;
		end

reg Pass_3;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_3<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1140==mem[3])&&(Pass_2))
				Pass_3<=1;
			else
				Pass_3<=0;
		end

reg Pass_4;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_4<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1150==mem[4])&&(Pass_3))
				Pass_4<=1;
			else
				Pass_4<=0;
		end

reg Pass_5;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_5<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1160==mem[5])&&(Pass_4))
				Pass_5<=1;
			else
				Pass_5<=0;
		end

reg Pass_6;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_6<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1170==mem[6])&&(Pass_5))
				Pass_6<=1;
			else
				Pass_6<=0;
		end

reg Pass_7;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_7<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1180==mem[7])&&(Pass_6))
				Pass_7<=1;
			else
				Pass_7<=0;
		end

reg Pass_8;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_8<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1190==mem[8])&&(Pass_7))
				Pass_8<=1;
			else
				Pass_8<=0;
		end

reg Pass_9;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_9<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11A0==mem[9])&&(Pass_8))
				Pass_9<=1;
			else
				Pass_9<=0;
		end

reg Pass_10;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_10<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11B0==mem[10])&&(Pass_9))
				Pass_10<=1;
			else
				Pass_10<=0;
		end

reg Pass_11;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_11<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11C0==mem[11])&&(Pass_10))
				Pass_11<=1;
			else
				Pass_11<=0;
		end

reg Pass_12;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_12<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11D0==mem[12])&&(Pass_11))
				Pass_12<=1;
			else
				Pass_12<=0;
		end

reg Pass_13;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_13<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11E0==mem[13])&&(Pass_12))
				Pass_13<=1;
			else
				Pass_13<=0;
		end

reg Pass_14;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_14<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1210==mem[14])&&(Pass_13))
				Pass_14<=1;
			else
				Pass_14<=0;
		end

reg Pass_15;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_15<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1220==mem[15])&&(Pass_14))
				Pass_15<=1;
			else
				Pass_15<=0;
		end

reg Pass_16;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_16<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1230==mem[16])&&(Pass_15))
				Pass_16<=1;
			else
				Pass_16<=0;
		end

reg Pass_17;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_17<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1240==mem[17])&&(Pass_16))
				Pass_17<=1;
			else
				Pass_17<=0;
		end

reg Pass_18;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_18<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1250==mem[18])&&(Pass_17))
				Pass_18<=1;
			else
				Pass_18<=0;
		end

reg Pass_19;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_19<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1260==mem[19])&&(Pass_18))
				Pass_19<=1;
			else
				Pass_19<=0;
		end

reg Pass_20;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_20<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1270==mem[20])&&(Pass_19))
				Pass_20<=1;
			else
				Pass_20<=0;
		end

reg Pass_21;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_21<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1280==mem[21])&&(Pass_20))
				Pass_21<=1;
			else
				Pass_21<=0;
		end

reg Pass_22;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_22<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1290==mem[22])&&(Pass_21))
				Pass_22<=1;
			else
				Pass_22<=0;
		end

reg Pass_23;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_23<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12A0==mem[23])&&(Pass_22))
				Pass_23<=1;
			else
				Pass_23<=0;
		end

reg Pass_24;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_24<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12B0==mem[24])&&(Pass_23))
				Pass_24<=1;
			else
				Pass_24<=0;
		end

reg Pass_25;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_25<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12C0==mem[25])&&(Pass_24))
				Pass_25<=1;
			else
				Pass_25<=0;
		end

reg Pass_26;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_26<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12D0==mem[26])&&(Pass_25))
				Pass_26<=1;
			else
				Pass_26<=0;
		end

reg Pass_27;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_27<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12E0==mem[27])&&(Pass_26))
				Pass_27<=1;
			else
				Pass_27<=0;
		end

reg Pass_28;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_28<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1310==mem[28])&&(Pass_27))
				Pass_28<=1;
			else
				Pass_28<=0;
		end

reg Pass_29;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_29<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1320==mem[29])&&(Pass_28))
				Pass_29<=1;
			else
				Pass_29<=0;
		end

reg Pass_30;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_30<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1330==mem[30])&&(Pass_29))
				Pass_30<=1;
			else
				Pass_30<=0;
		end

reg Pass_31;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_31<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1340==mem[31])&&(Pass_30))
				Pass_31<=1;
			else
				Pass_31<=0;
		end

reg Pass_32;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_32<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1350==mem[32])&&(Pass_31))
				Pass_32<=1;
			else
				Pass_32<=0;
		end

reg Pass_33;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_33<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1360==mem[33])&&(Pass_32))
				Pass_33<=1;
			else
				Pass_33<=0;
		end

reg Pass_34;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_34<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1370==mem[34])&&(Pass_33))
				Pass_34<=1;
			else
				Pass_34<=0;
		end

reg Pass_35;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_35<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1380==mem[35])&&(Pass_34))
				Pass_35<=1;
			else
				Pass_35<=0;
		end

reg Pass_36;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_36<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1390==mem[36])&&(Pass_35))
				Pass_36<=1;
			else
				Pass_36<=0;
		end

reg Pass_37;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_37<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13A0==mem[37])&&(Pass_36))
				Pass_37<=1;
			else
				Pass_37<=0;
		end

reg Pass_38;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_38<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13B0==mem[38])&&(Pass_37))
				Pass_38<=1;
			else
				Pass_38<=0;
		end

reg Pass_39;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_39<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13C0==mem[39])&&(Pass_38))
				Pass_39<=1;
			else
				Pass_39<=0;
		end

reg Pass_40;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_40<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13D0==mem[40])&&(Pass_39))
				Pass_40<=1;
			else
				Pass_40<=0;
		end

reg Pass_41;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_41<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13E0==mem[41])&&(Pass_40))
				Pass_41<=1;
			else
				Pass_41<=0;
		end

reg Pass_42;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_42<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1410==mem[42])&&(Pass_41))
				Pass_42<=1;
			else
				Pass_42<=0;
		end

reg Pass_43;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_43<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1420==mem[43])&&(Pass_42))
				Pass_43<=1;
			else
				Pass_43<=0;
		end

reg Pass_44;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_44<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1430==mem[44])&&(Pass_43))
				Pass_44<=1;
			else
				Pass_44<=0;
		end

reg Pass_45;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_45<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1440==mem[45])&&(Pass_44))
				Pass_45<=1;
			else
				Pass_45<=0;
		end

reg Pass_46;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_46<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1450==mem[46])&&(Pass_45))
				Pass_46<=1;
			else
				Pass_46<=0;
		end

reg Pass_47;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_47<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1460==mem[47])&&(Pass_46))
				Pass_47<=1;
			else
				Pass_47<=0;
		end

reg Pass_48;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_48<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1470==mem[48])&&(Pass_47))
				Pass_48<=1;
			else
				Pass_48<=0;
		end

reg Pass_49;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_49<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1480==mem[49])&&(Pass_48))
				Pass_49<=1;
			else
				Pass_49<=0;
		end

reg Pass_50;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_50<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1490==mem[50])&&(Pass_49))
				Pass_50<=1;
			else
				Pass_50<=0;
		end

reg Pass_51;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_51<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14A0==mem[51])&&(Pass_50))
				Pass_51<=1;
			else
				Pass_51<=0;
		end

reg Pass_52;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_52<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14B0==mem[52])&&(Pass_51))
				Pass_52<=1;
			else
				Pass_52<=0;
		end

reg Pass_53;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_53<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14C0==mem[53])&&(Pass_52))
				Pass_53<=1;
			else
				Pass_53<=0;
		end

reg Pass_54;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_54<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14D0==mem[54])&&(Pass_53))
				Pass_54<=1;
			else
				Pass_54<=0;
		end

reg Pass_55;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_55<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14E0==mem[55])&&(Pass_54))
				Pass_55<=1;
			else
				Pass_55<=0;
		end

reg Pass_56;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_56<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1510==mem[56])&&(Pass_55))
				Pass_56<=1;
			else
				Pass_56<=0;
		end

reg Pass_57;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_57<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1520==mem[57])&&(Pass_56))
				Pass_57<=1;
			else
				Pass_57<=0;
		end

reg Pass_58;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_58<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1530==mem[58])&&(Pass_57))
				Pass_58<=1;
			else
				Pass_58<=0;
		end

reg Pass_59;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_59<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1540==mem[59])&&(Pass_58))
				Pass_59<=1;
			else
				Pass_59<=0;
		end

reg Pass_60;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_60<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1550==mem[60])&&(Pass_59))
				Pass_60<=1;
			else
				Pass_60<=0;
		end

reg Pass_61;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_61<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1560==mem[61])&&(Pass_60))
				Pass_61<=1;
			else
				Pass_61<=0;
		end

reg Pass_62;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_62<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1570==mem[62])&&(Pass_61))
				Pass_62<=1;
			else
				Pass_62<=0;
		end

reg Pass_63;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_63<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1580==mem[63])&&(Pass_62))
				Pass_63<=1;
			else
				Pass_63<=0;
		end

reg Pass_64;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_64<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1590==mem[64])&&(Pass_63))
				Pass_64<=1;
			else
				Pass_64<=0;
		end

reg Pass_65;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_65<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15A0==mem[65])&&(Pass_64))
				Pass_65<=1;
			else
				Pass_65<=0;
		end

reg Pass_66;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_66<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15B0==mem[66])&&(Pass_65))
				Pass_66<=1;
			else
				Pass_66<=0;
		end

reg Pass_67;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_67<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15C0==mem[67])&&(Pass_66))
				Pass_67<=1;
			else
				Pass_67<=0;
		end

reg Pass_68;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_68<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15D0==mem[68])&&(Pass_67))
				Pass_68<=1;
			else
				Pass_68<=0;
		end

reg Pass_69;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_69<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15E0==mem[69])&&(Pass_68))
				Pass_69<=1;
			else
				Pass_69<=0;
		end

reg Pass_70;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_70<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1610==mem[70])&&(Pass_69))
				Pass_70<=1;
			else
				Pass_70<=0;
		end

reg Pass_71;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_71<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1620==mem[71])&&(Pass_70))
				Pass_71<=1;
			else
				Pass_71<=0;
		end

reg Pass_72;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_72<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1630==mem[72])&&(Pass_71))
				Pass_72<=1;
			else
				Pass_72<=0;
		end

reg Pass_73;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_73<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1640==mem[73])&&(Pass_72))
				Pass_73<=1;
			else
				Pass_73<=0;
		end

reg Pass_74;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_74<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1650==mem[74])&&(Pass_73))
				Pass_74<=1;
			else
				Pass_74<=0;
		end

reg Pass_75;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_75<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1660==mem[75])&&(Pass_74))
				Pass_75<=1;
			else
				Pass_75<=0;
		end

reg Pass_76;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_76<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1670==mem[76])&&(Pass_75))
				Pass_76<=1;
			else
				Pass_76<=0;
		end

reg Pass_77;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_77<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1680==mem[77])&&(Pass_76))
				Pass_77<=1;
			else
				Pass_77<=0;
		end

reg Pass_78;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_78<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1690==mem[78])&&(Pass_77))
				Pass_78<=1;
			else
				Pass_78<=0;
		end

reg Pass_79;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_79<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16A0==mem[79])&&(Pass_78))
				Pass_79<=1;
			else
				Pass_79<=0;
		end

reg Pass_80;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_80<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16B0==mem[80])&&(Pass_79))
				Pass_80<=1;
			else
				Pass_80<=0;
		end

reg Pass_81;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_81<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16C0==mem[81])&&(Pass_80))
				Pass_81<=1;
			else
				Pass_81<=0;
		end

reg Pass_82;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_82<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16D0==mem[82])&&(Pass_81))
				Pass_82<=1;
			else
				Pass_82<=0;
		end

reg Pass_83;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_83<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16E0==mem[83])&&(Pass_82))
				Pass_83<=1;
			else
				Pass_83<=0;
		end

reg Pass_84;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_84<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1710==mem[84])&&(Pass_83))
				Pass_84<=1;
			else
				Pass_84<=0;
		end

reg Pass_85;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_85<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1720==mem[85])&&(Pass_84))
				Pass_85<=1;
			else
				Pass_85<=0;
		end

reg Pass_86;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_86<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1730==mem[86])&&(Pass_85))
				Pass_86<=1;
			else
				Pass_86<=0;
		end

reg Pass_87;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_87<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1740==mem[87])&&(Pass_86))
				Pass_87<=1;
			else
				Pass_87<=0;
		end

reg Pass_88;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_88<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1750==mem[88])&&(Pass_87))
				Pass_88<=1;
			else
				Pass_88<=0;
		end

reg Pass_89;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_89<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1760==mem[89])&&(Pass_88))
				Pass_89<=1;
			else
				Pass_89<=0;
		end

reg Pass_90;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_90<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1770==mem[90])&&(Pass_89))
				Pass_90<=1;
			else
				Pass_90<=0;
		end

reg Pass_91;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_91<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1780==mem[91])&&(Pass_90))
				Pass_91<=1;
			else
				Pass_91<=0;
		end

reg Pass_92;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_92<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1790==mem[92])&&(Pass_91))
				Pass_92<=1;
			else
				Pass_92<=0;
		end

reg Pass_93;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_93<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17A0==mem[93])&&(Pass_92))
				Pass_93<=1;
			else
				Pass_93<=0;
		end

reg Pass_94;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_94<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17B0==mem[94])&&(Pass_93))
				Pass_94<=1;
			else
				Pass_94<=0;
		end

reg Pass_95;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_95<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17C0==mem[95])&&(Pass_94))
				Pass_95<=1;
			else
				Pass_95<=0;
		end

reg Pass_96;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_96<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17D0==mem[96])&&(Pass_95))
				Pass_96<=1;
			else
				Pass_96<=0;
		end

reg Pass_97;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_97<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17E0==mem[97])&&(Pass_96))
				Pass_97<=1;
			else
				Pass_97<=0;
		end

reg Pass_98;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_98<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1810==mem[98])&&(Pass_97))
				Pass_98<=1;
			else
				Pass_98<=0;
		end

reg Pass_99;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_99<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1820==mem[99])&&(Pass_98))
				Pass_99<=1;
			else
				Pass_99<=0;
		end

reg Pass_100;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_100<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1830==mem[100])&&(Pass_99))
				Pass_100<=1;
			else
				Pass_100<=0;
		end

reg Pass_101;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_101<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1840==mem[101])&&(Pass_100))
				Pass_101<=1;
			else
				Pass_101<=0;
		end

reg Pass_102;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_102<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1850==mem[102])&&(Pass_101))
				Pass_102<=1;
			else
				Pass_102<=0;
		end

reg Pass_103;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_103<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1860==mem[103])&&(Pass_102))
				Pass_103<=1;
			else
				Pass_103<=0;
		end

reg Pass_104;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_104<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1870==mem[104])&&(Pass_103))
				Pass_104<=1;
			else
				Pass_104<=0;
		end

reg Pass_105;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_105<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1880==mem[105])&&(Pass_104))
				Pass_105<=1;
			else
				Pass_105<=0;
		end

reg Pass_106;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_106<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1890==mem[106])&&(Pass_105))
				Pass_106<=1;
			else
				Pass_106<=0;
		end

reg Pass_107;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_107<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18A0==mem[107])&&(Pass_106))
				Pass_107<=1;
			else
				Pass_107<=0;
		end

reg Pass_108;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_108<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18B0==mem[108])&&(Pass_107))
				Pass_108<=1;
			else
				Pass_108<=0;
		end

reg Pass_109;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_109<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18C0==mem[109])&&(Pass_108))
				Pass_109<=1;
			else
				Pass_109<=0;
		end

reg Pass_110;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_110<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18D0==mem[110])&&(Pass_109))
				Pass_110<=1;
			else
				Pass_110<=0;
		end

reg Pass_111;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_111<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18E0==mem[111])&&(Pass_110))
				Pass_111<=1;
			else
				Pass_111<=0;
		end

reg Pass_112;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_112<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1910==mem[112])&&(Pass_111))
				Pass_112<=1;
			else
				Pass_112<=0;
		end

reg Pass_113;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_113<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1920==mem[113])&&(Pass_112))
				Pass_113<=1;
			else
				Pass_113<=0;
		end

reg Pass_114;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_114<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1930==mem[114])&&(Pass_113))
				Pass_114<=1;
			else
				Pass_114<=0;
		end

reg Pass_115;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_115<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1940==mem[115])&&(Pass_114))
				Pass_115<=1;
			else
				Pass_115<=0;
		end

reg Pass_116;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_116<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1950==mem[116])&&(Pass_115))
				Pass_116<=1;
			else
				Pass_116<=0;
		end

reg Pass_117;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_117<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1960==mem[117])&&(Pass_116))
				Pass_117<=1;
			else
				Pass_117<=0;
		end

reg Pass_118;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_118<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1970==mem[118])&&(Pass_117))
				Pass_118<=1;
			else
				Pass_118<=0;
		end

reg Pass_119;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_119<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1980==mem[119])&&(Pass_118))
				Pass_119<=1;
			else
				Pass_119<=0;
		end

reg Pass_120;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_120<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1990==mem[120])&&(Pass_119))
				Pass_120<=1;
			else
				Pass_120<=0;
		end

reg Pass_121;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_121<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19A0==mem[121])&&(Pass_120))
				Pass_121<=1;
			else
				Pass_121<=0;
		end

reg Pass_122;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_122<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19B0==mem[122])&&(Pass_121))
				Pass_122<=1;
			else
				Pass_122<=0;
		end

reg Pass_123;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_123<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19C0==mem[123])&&(Pass_122))
				Pass_123<=1;
			else
				Pass_123<=0;
		end

reg Pass_124;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_124<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19D0==mem[124])&&(Pass_123))
				Pass_124<=1;
			else
				Pass_124<=0;
		end

reg Pass_125;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_125<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19E0==mem[125])&&(Pass_124))
				Pass_125<=1;
			else
				Pass_125<=0;
		end

reg Pass_126;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_126<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A10==mem[126])&&(Pass_125))
				Pass_126<=1;
			else
				Pass_126<=0;
		end

reg Pass_127;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_127<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A20==mem[127])&&(Pass_126))
				Pass_127<=1;
			else
				Pass_127<=0;
		end

reg Pass_128;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_128<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A30==mem[128])&&(Pass_127))
				Pass_128<=1;
			else
				Pass_128<=0;
		end

reg Pass_129;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_129<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A40==mem[129])&&(Pass_128))
				Pass_129<=1;
			else
				Pass_129<=0;
		end

reg Pass_130;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_130<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A50==mem[130])&&(Pass_129))
				Pass_130<=1;
			else
				Pass_130<=0;
		end

reg Pass_131;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_131<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A60==mem[131])&&(Pass_130))
				Pass_131<=1;
			else
				Pass_131<=0;
		end

reg Pass_132;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_132<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A70==mem[132])&&(Pass_131))
				Pass_132<=1;
			else
				Pass_132<=0;
		end

reg Pass_133;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_133<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A80==mem[133])&&(Pass_132))
				Pass_133<=1;
			else
				Pass_133<=0;
		end

reg Pass_134;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_134<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A90==mem[134])&&(Pass_133))
				Pass_134<=1;
			else
				Pass_134<=0;
		end

reg Pass_135;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_135<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AA0==mem[135])&&(Pass_134))
				Pass_135<=1;
			else
				Pass_135<=0;
		end

reg Pass_136;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_136<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AB0==mem[136])&&(Pass_135))
				Pass_136<=1;
			else
				Pass_136<=0;
		end

reg Pass_137;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_137<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AC0==mem[137])&&(Pass_136))
				Pass_137<=1;
			else
				Pass_137<=0;
		end

reg Pass_138;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_138<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AD0==mem[138])&&(Pass_137))
				Pass_138<=1;
			else
				Pass_138<=0;
		end

reg Pass_139;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_139<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AE0==mem[139])&&(Pass_138))
				Pass_139<=1;
			else
				Pass_139<=0;
		end

reg Pass_140;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_140<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B10==mem[140])&&(Pass_139))
				Pass_140<=1;
			else
				Pass_140<=0;
		end

reg Pass_141;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_141<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B20==mem[141])&&(Pass_140))
				Pass_141<=1;
			else
				Pass_141<=0;
		end

reg Pass_142;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_142<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B30==mem[142])&&(Pass_141))
				Pass_142<=1;
			else
				Pass_142<=0;
		end

reg Pass_143;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_143<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B40==mem[143])&&(Pass_142))
				Pass_143<=1;
			else
				Pass_143<=0;
		end

reg Pass_144;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_144<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B50==mem[144])&&(Pass_143))
				Pass_144<=1;
			else
				Pass_144<=0;
		end

reg Pass_145;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_145<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B60==mem[145])&&(Pass_144))
				Pass_145<=1;
			else
				Pass_145<=0;
		end

reg Pass_146;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_146<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B70==mem[146])&&(Pass_145))
				Pass_146<=1;
			else
				Pass_146<=0;
		end

reg Pass_147;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_147<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B80==mem[147])&&(Pass_146))
				Pass_147<=1;
			else
				Pass_147<=0;
		end

reg Pass_148;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_148<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B90==mem[148])&&(Pass_147))
				Pass_148<=1;
			else
				Pass_148<=0;
		end

reg Pass_149;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_149<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BA0==mem[149])&&(Pass_148))
				Pass_149<=1;
			else
				Pass_149<=0;
		end

reg Pass_150;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_150<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BB0==mem[150])&&(Pass_149))
				Pass_150<=1;
			else
				Pass_150<=0;
		end

reg Pass_151;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_151<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BC0==mem[151])&&(Pass_150))
				Pass_151<=1;
			else
				Pass_151<=0;
		end

reg Pass_152;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_152<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BD0==mem[152])&&(Pass_151))
				Pass_152<=1;
			else
				Pass_152<=0;
		end

reg Pass_153;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_153<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BE0==mem[153])&&(Pass_152))
				Pass_153<=1;
			else
				Pass_153<=0;
		end

reg Pass_154;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_154<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C10==mem[154])&&(Pass_153))
				Pass_154<=1;
			else
				Pass_154<=0;
		end

reg Pass_155;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_155<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C20==mem[155])&&(Pass_154))
				Pass_155<=1;
			else
				Pass_155<=0;
		end

reg Pass_156;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_156<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C30==mem[156])&&(Pass_155))
				Pass_156<=1;
			else
				Pass_156<=0;
		end

reg Pass_157;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_157<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C40==mem[157])&&(Pass_156))
				Pass_157<=1;
			else
				Pass_157<=0;
		end

reg Pass_158;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_158<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C50==mem[158])&&(Pass_157))
				Pass_158<=1;
			else
				Pass_158<=0;
		end

reg Pass_159;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_159<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C60==mem[159])&&(Pass_158))
				Pass_159<=1;
			else
				Pass_159<=0;
		end

reg Pass_160;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_160<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C70==mem[160])&&(Pass_159))
				Pass_160<=1;
			else
				Pass_160<=0;
		end

reg Pass_161;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_161<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C80==mem[161])&&(Pass_160))
				Pass_161<=1;
			else
				Pass_161<=0;
		end

reg Pass_162;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_162<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C90==mem[162])&&(Pass_161))
				Pass_162<=1;
			else
				Pass_162<=0;
		end

reg Pass_163;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_163<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CA0==mem[163])&&(Pass_162))
				Pass_163<=1;
			else
				Pass_163<=0;
		end

reg Pass_164;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_164<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CB0==mem[164])&&(Pass_163))
				Pass_164<=1;
			else
				Pass_164<=0;
		end

reg Pass_165;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_165<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CC0==mem[165])&&(Pass_164))
				Pass_165<=1;
			else
				Pass_165<=0;
		end

reg Pass_166;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_166<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CD0==mem[166])&&(Pass_165))
				Pass_166<=1;
			else
				Pass_166<=0;
		end

reg Pass_167;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_167<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CE0==mem[167])&&(Pass_166))
				Pass_167<=1;
			else
				Pass_167<=0;
		end

reg Pass_168;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_168<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D10==mem[168])&&(Pass_167))
				Pass_168<=1;
			else
				Pass_168<=0;
		end

reg Pass_169;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_169<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D20==mem[169])&&(Pass_168))
				Pass_169<=1;
			else
				Pass_169<=0;
		end

reg Pass_170;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_170<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D30==mem[170])&&(Pass_169))
				Pass_170<=1;
			else
				Pass_170<=0;
		end

reg Pass_171;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_171<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D40==mem[171])&&(Pass_170))
				Pass_171<=1;
			else
				Pass_171<=0;
		end

reg Pass_172;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_172<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D50==mem[172])&&(Pass_171))
				Pass_172<=1;
			else
				Pass_172<=0;
		end

reg Pass_173;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_173<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D60==mem[173])&&(Pass_172))
				Pass_173<=1;
			else
				Pass_173<=0;
		end

reg Pass_174;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_174<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D70==mem[174])&&(Pass_173))
				Pass_174<=1;
			else
				Pass_174<=0;
		end

reg Pass_175;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_175<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D80==mem[175])&&(Pass_174))
				Pass_175<=1;
			else
				Pass_175<=0;
		end

reg Pass_176;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_176<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D90==mem[176])&&(Pass_175))
				Pass_176<=1;
			else
				Pass_176<=0;
		end

reg Pass_177;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_177<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DA0==mem[177])&&(Pass_176))
				Pass_177<=1;
			else
				Pass_177<=0;
		end

reg Pass_178;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_178<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DB0==mem[178])&&(Pass_177))
				Pass_178<=1;
			else
				Pass_178<=0;
		end

reg Pass_179;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_179<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DC0==mem[179])&&(Pass_178))
				Pass_179<=1;
			else
				Pass_179<=0;
		end

reg Pass_180;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_180<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DD0==mem[180])&&(Pass_179))
				Pass_180<=1;
			else
				Pass_180<=0;
		end

reg Pass_181;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_181<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DE0==mem[181])&&(Pass_180))
				Pass_181<=1;
			else
				Pass_181<=0;
		end

reg Pass_182;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_182<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E10==mem[182])&&(Pass_181))
				Pass_182<=1;
			else
				Pass_182<=0;
		end

reg Pass_183;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_183<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E20==mem[183])&&(Pass_182))
				Pass_183<=1;
			else
				Pass_183<=0;
		end

reg Pass_184;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_184<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E30==mem[184])&&(Pass_183))
				Pass_184<=1;
			else
				Pass_184<=0;
		end

reg Pass_185;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_185<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E40==mem[185])&&(Pass_184))
				Pass_185<=1;
			else
				Pass_185<=0;
		end

reg Pass_186;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_186<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E50==mem[186])&&(Pass_185))
				Pass_186<=1;
			else
				Pass_186<=0;
		end

reg Pass_187;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_187<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E60==mem[187])&&(Pass_186))
				Pass_187<=1;
			else
				Pass_187<=0;
		end

reg Pass_188;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_188<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E70==mem[188])&&(Pass_187))
				Pass_188<=1;
			else
				Pass_188<=0;
		end

reg Pass_189;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_189<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E80==mem[189])&&(Pass_188))
				Pass_189<=1;
			else
				Pass_189<=0;
		end

reg Pass_190;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_190<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E90==mem[190])&&(Pass_189))
				Pass_190<=1;
			else
				Pass_190<=0;
		end

reg Pass_191;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_191<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1EA0==mem[191])&&(Pass_190))
				Pass_191<=1;
			else
				Pass_191<=0;
		end

reg Pass_192;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_192<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1EB0==mem[192])&&(Pass_191))
				Pass_192<=1;
			else
				Pass_192<=0;
		end

reg Pass_193;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_193<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1EC0==mem[193])&&(Pass_192))
				Pass_193<=1;
			else
				Pass_193<=0;
		end

reg Pass_194;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_194<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1ED0==mem[194])&&(Pass_193))
				Pass_194<=1;
			else
				Pass_194<=0;
		end

reg Pass_195;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_195<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1EE0==mem[195])&&(Pass_194))
				Pass_195<=1;
			else
				Pass_195<=0;
		end

reg Pass_196;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_196<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1111==mem[196])&&(Pass_195))
				Pass_196<=1;
			else
				Pass_196<=0;
		end

reg Pass_197;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_197<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1121==mem[197])&&(Pass_196))
				Pass_197<=1;
			else
				Pass_197<=0;
		end

reg Pass_198;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_198<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1131==mem[198])&&(Pass_197))
				Pass_198<=1;
			else
				Pass_198<=0;
		end

reg Pass_199;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_199<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1141==mem[199])&&(Pass_198))
				Pass_199<=1;
			else
				Pass_199<=0;
		end

reg Pass_200;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_200<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1151==mem[200])&&(Pass_199))
				Pass_200<=1;
			else
				Pass_200<=0;
		end

reg Pass_201;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_201<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1161==mem[201])&&(Pass_200))
				Pass_201<=1;
			else
				Pass_201<=0;
		end

reg Pass_202;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_202<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1171==mem[202])&&(Pass_201))
				Pass_202<=1;
			else
				Pass_202<=0;
		end

reg Pass_203;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_203<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1181==mem[203])&&(Pass_202))
				Pass_203<=1;
			else
				Pass_203<=0;
		end

reg Pass_204;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_204<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1191==mem[204])&&(Pass_203))
				Pass_204<=1;
			else
				Pass_204<=0;
		end

reg Pass_205;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_205<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11A1==mem[205])&&(Pass_204))
				Pass_205<=1;
			else
				Pass_205<=0;
		end

reg Pass_206;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_206<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11B1==mem[206])&&(Pass_205))
				Pass_206<=1;
			else
				Pass_206<=0;
		end

reg Pass_207;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_207<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11C1==mem[207])&&(Pass_206))
				Pass_207<=1;
			else
				Pass_207<=0;
		end

reg Pass_208;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_208<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11D1==mem[208])&&(Pass_207))
				Pass_208<=1;
			else
				Pass_208<=0;
		end

reg Pass_209;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_209<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11E1==mem[209])&&(Pass_208))
				Pass_209<=1;
			else
				Pass_209<=0;
		end

reg Pass_210;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_210<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1211==mem[210])&&(Pass_209))
				Pass_210<=1;
			else
				Pass_210<=0;
		end

reg Pass_211;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_211<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1221==mem[211])&&(Pass_210))
				Pass_211<=1;
			else
				Pass_211<=0;
		end

reg Pass_212;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_212<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1231==mem[212])&&(Pass_211))
				Pass_212<=1;
			else
				Pass_212<=0;
		end

reg Pass_213;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_213<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1241==mem[213])&&(Pass_212))
				Pass_213<=1;
			else
				Pass_213<=0;
		end

reg Pass_214;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_214<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1251==mem[214])&&(Pass_213))
				Pass_214<=1;
			else
				Pass_214<=0;
		end

reg Pass_215;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_215<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1261==mem[215])&&(Pass_214))
				Pass_215<=1;
			else
				Pass_215<=0;
		end

reg Pass_216;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_216<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1271==mem[216])&&(Pass_215))
				Pass_216<=1;
			else
				Pass_216<=0;
		end

reg Pass_217;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_217<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1281==mem[217])&&(Pass_216))
				Pass_217<=1;
			else
				Pass_217<=0;
		end

reg Pass_218;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_218<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1291==mem[218])&&(Pass_217))
				Pass_218<=1;
			else
				Pass_218<=0;
		end

reg Pass_219;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_219<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12A1==mem[219])&&(Pass_218))
				Pass_219<=1;
			else
				Pass_219<=0;
		end

reg Pass_220;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_220<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12B1==mem[220])&&(Pass_219))
				Pass_220<=1;
			else
				Pass_220<=0;
		end

reg Pass_221;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_221<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12C1==mem[221])&&(Pass_220))
				Pass_221<=1;
			else
				Pass_221<=0;
		end

reg Pass_222;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_222<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12D1==mem[222])&&(Pass_221))
				Pass_222<=1;
			else
				Pass_222<=0;
		end

reg Pass_223;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_223<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12E1==mem[223])&&(Pass_222))
				Pass_223<=1;
			else
				Pass_223<=0;
		end

reg Pass_224;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_224<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1311==mem[224])&&(Pass_223))
				Pass_224<=1;
			else
				Pass_224<=0;
		end

reg Pass_225;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_225<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1321==mem[225])&&(Pass_224))
				Pass_225<=1;
			else
				Pass_225<=0;
		end

reg Pass_226;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_226<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1331==mem[226])&&(Pass_225))
				Pass_226<=1;
			else
				Pass_226<=0;
		end

reg Pass_227;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_227<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1341==mem[227])&&(Pass_226))
				Pass_227<=1;
			else
				Pass_227<=0;
		end

reg Pass_228;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_228<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1351==mem[228])&&(Pass_227))
				Pass_228<=1;
			else
				Pass_228<=0;
		end

reg Pass_229;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_229<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1361==mem[229])&&(Pass_228))
				Pass_229<=1;
			else
				Pass_229<=0;
		end

reg Pass_230;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_230<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1371==mem[230])&&(Pass_229))
				Pass_230<=1;
			else
				Pass_230<=0;
		end

reg Pass_231;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_231<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1381==mem[231])&&(Pass_230))
				Pass_231<=1;
			else
				Pass_231<=0;
		end

reg Pass_232;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_232<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1391==mem[232])&&(Pass_231))
				Pass_232<=1;
			else
				Pass_232<=0;
		end

reg Pass_233;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_233<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13A1==mem[233])&&(Pass_232))
				Pass_233<=1;
			else
				Pass_233<=0;
		end

reg Pass_234;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_234<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13B1==mem[234])&&(Pass_233))
				Pass_234<=1;
			else
				Pass_234<=0;
		end

reg Pass_235;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_235<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13C1==mem[235])&&(Pass_234))
				Pass_235<=1;
			else
				Pass_235<=0;
		end

reg Pass_236;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_236<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13D1==mem[236])&&(Pass_235))
				Pass_236<=1;
			else
				Pass_236<=0;
		end

reg Pass_237;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_237<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13E1==mem[237])&&(Pass_236))
				Pass_237<=1;
			else
				Pass_237<=0;
		end

reg Pass_238;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_238<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1411==mem[238])&&(Pass_237))
				Pass_238<=1;
			else
				Pass_238<=0;
		end

reg Pass_239;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_239<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1421==mem[239])&&(Pass_238))
				Pass_239<=1;
			else
				Pass_239<=0;
		end

reg Pass_240;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_240<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1431==mem[240])&&(Pass_239))
				Pass_240<=1;
			else
				Pass_240<=0;
		end

reg Pass_241;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_241<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1441==mem[241])&&(Pass_240))
				Pass_241<=1;
			else
				Pass_241<=0;
		end

reg Pass_242;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_242<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1451==mem[242])&&(Pass_241))
				Pass_242<=1;
			else
				Pass_242<=0;
		end

reg Pass_243;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_243<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1461==mem[243])&&(Pass_242))
				Pass_243<=1;
			else
				Pass_243<=0;
		end

reg Pass_244;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_244<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1471==mem[244])&&(Pass_243))
				Pass_244<=1;
			else
				Pass_244<=0;
		end

reg Pass_245;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_245<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1481==mem[245])&&(Pass_244))
				Pass_245<=1;
			else
				Pass_245<=0;
		end

reg Pass_246;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_246<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1491==mem[246])&&(Pass_245))
				Pass_246<=1;
			else
				Pass_246<=0;
		end

reg Pass_247;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_247<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14A1==mem[247])&&(Pass_246))
				Pass_247<=1;
			else
				Pass_247<=0;
		end

reg Pass_248;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_248<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14B1==mem[248])&&(Pass_247))
				Pass_248<=1;
			else
				Pass_248<=0;
		end

reg Pass_249;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_249<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14C1==mem[249])&&(Pass_248))
				Pass_249<=1;
			else
				Pass_249<=0;
		end

reg Pass_250;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_250<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14D1==mem[250])&&(Pass_249))
				Pass_250<=1;
			else
				Pass_250<=0;
		end

reg Pass_251;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_251<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14E1==mem[251])&&(Pass_250))
				Pass_251<=1;
			else
				Pass_251<=0;
		end

reg Pass_252;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_252<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1511==mem[252])&&(Pass_251))
				Pass_252<=1;
			else
				Pass_252<=0;
		end

reg Pass_253;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_253<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1521==mem[253])&&(Pass_252))
				Pass_253<=1;
			else
				Pass_253<=0;
		end

reg Pass_254;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_254<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1531==mem[254])&&(Pass_253))
				Pass_254<=1;
			else
				Pass_254<=0;
		end

reg Pass_255;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_255<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1541==mem[255])&&(Pass_254))
				Pass_255<=1;
			else
				Pass_255<=0;
		end

reg Pass_256;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_256<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1551==mem[256])&&(Pass_255))
				Pass_256<=1;
			else
				Pass_256<=0;
		end

reg Pass_257;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_257<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1561==mem[257])&&(Pass_256))
				Pass_257<=1;
			else
				Pass_257<=0;
		end

reg Pass_258;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_258<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1571==mem[258])&&(Pass_257))
				Pass_258<=1;
			else
				Pass_258<=0;
		end

reg Pass_259;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_259<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1581==mem[259])&&(Pass_258))
				Pass_259<=1;
			else
				Pass_259<=0;
		end

reg Pass_260;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_260<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1591==mem[260])&&(Pass_259))
				Pass_260<=1;
			else
				Pass_260<=0;
		end

reg Pass_261;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_261<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15A1==mem[261])&&(Pass_260))
				Pass_261<=1;
			else
				Pass_261<=0;
		end

reg Pass_262;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_262<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15B1==mem[262])&&(Pass_261))
				Pass_262<=1;
			else
				Pass_262<=0;
		end

reg Pass_263;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_263<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15C1==mem[263])&&(Pass_262))
				Pass_263<=1;
			else
				Pass_263<=0;
		end

reg Pass_264;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_264<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15D1==mem[264])&&(Pass_263))
				Pass_264<=1;
			else
				Pass_264<=0;
		end

reg Pass_265;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_265<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15E1==mem[265])&&(Pass_264))
				Pass_265<=1;
			else
				Pass_265<=0;
		end

reg Pass_266;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_266<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1611==mem[266])&&(Pass_265))
				Pass_266<=1;
			else
				Pass_266<=0;
		end

reg Pass_267;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_267<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1621==mem[267])&&(Pass_266))
				Pass_267<=1;
			else
				Pass_267<=0;
		end

reg Pass_268;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_268<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1631==mem[268])&&(Pass_267))
				Pass_268<=1;
			else
				Pass_268<=0;
		end

reg Pass_269;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_269<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1641==mem[269])&&(Pass_268))
				Pass_269<=1;
			else
				Pass_269<=0;
		end

reg Pass_270;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_270<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1651==mem[270])&&(Pass_269))
				Pass_270<=1;
			else
				Pass_270<=0;
		end

reg Pass_271;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_271<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1661==mem[271])&&(Pass_270))
				Pass_271<=1;
			else
				Pass_271<=0;
		end

reg Pass_272;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_272<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1671==mem[272])&&(Pass_271))
				Pass_272<=1;
			else
				Pass_272<=0;
		end

reg Pass_273;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_273<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1681==mem[273])&&(Pass_272))
				Pass_273<=1;
			else
				Pass_273<=0;
		end

reg Pass_274;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_274<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1691==mem[274])&&(Pass_273))
				Pass_274<=1;
			else
				Pass_274<=0;
		end

reg Pass_275;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_275<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16A1==mem[275])&&(Pass_274))
				Pass_275<=1;
			else
				Pass_275<=0;
		end

reg Pass_276;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_276<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16B1==mem[276])&&(Pass_275))
				Pass_276<=1;
			else
				Pass_276<=0;
		end

reg Pass_277;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_277<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16C1==mem[277])&&(Pass_276))
				Pass_277<=1;
			else
				Pass_277<=0;
		end

reg Pass_278;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_278<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16D1==mem[278])&&(Pass_277))
				Pass_278<=1;
			else
				Pass_278<=0;
		end

reg Pass_279;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_279<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16E1==mem[279])&&(Pass_278))
				Pass_279<=1;
			else
				Pass_279<=0;
		end

reg Pass_280;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_280<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1711==mem[280])&&(Pass_279))
				Pass_280<=1;
			else
				Pass_280<=0;
		end

reg Pass_281;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_281<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1721==mem[281])&&(Pass_280))
				Pass_281<=1;
			else
				Pass_281<=0;
		end

reg Pass_282;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_282<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1731==mem[282])&&(Pass_281))
				Pass_282<=1;
			else
				Pass_282<=0;
		end

reg Pass_283;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_283<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1741==mem[283])&&(Pass_282))
				Pass_283<=1;
			else
				Pass_283<=0;
		end

reg Pass_284;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_284<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1751==mem[284])&&(Pass_283))
				Pass_284<=1;
			else
				Pass_284<=0;
		end

reg Pass_285;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_285<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1761==mem[285])&&(Pass_284))
				Pass_285<=1;
			else
				Pass_285<=0;
		end

reg Pass_286;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_286<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1771==mem[286])&&(Pass_285))
				Pass_286<=1;
			else
				Pass_286<=0;
		end

reg Pass_287;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_287<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1781==mem[287])&&(Pass_286))
				Pass_287<=1;
			else
				Pass_287<=0;
		end

reg Pass_288;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_288<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1791==mem[288])&&(Pass_287))
				Pass_288<=1;
			else
				Pass_288<=0;
		end

reg Pass_289;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_289<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17A1==mem[289])&&(Pass_288))
				Pass_289<=1;
			else
				Pass_289<=0;
		end

reg Pass_290;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_290<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17B1==mem[290])&&(Pass_289))
				Pass_290<=1;
			else
				Pass_290<=0;
		end

reg Pass_291;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_291<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17C1==mem[291])&&(Pass_290))
				Pass_291<=1;
			else
				Pass_291<=0;
		end

reg Pass_292;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_292<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17D1==mem[292])&&(Pass_291))
				Pass_292<=1;
			else
				Pass_292<=0;
		end

reg Pass_293;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_293<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17E1==mem[293])&&(Pass_292))
				Pass_293<=1;
			else
				Pass_293<=0;
		end

reg Pass_294;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_294<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1811==mem[294])&&(Pass_293))
				Pass_294<=1;
			else
				Pass_294<=0;
		end

reg Pass_295;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_295<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1821==mem[295])&&(Pass_294))
				Pass_295<=1;
			else
				Pass_295<=0;
		end

reg Pass_296;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_296<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1831==mem[296])&&(Pass_295))
				Pass_296<=1;
			else
				Pass_296<=0;
		end

reg Pass_297;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_297<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1841==mem[297])&&(Pass_296))
				Pass_297<=1;
			else
				Pass_297<=0;
		end

reg Pass_298;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_298<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1851==mem[298])&&(Pass_297))
				Pass_298<=1;
			else
				Pass_298<=0;
		end

reg Pass_299;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_299<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1861==mem[299])&&(Pass_298))
				Pass_299<=1;
			else
				Pass_299<=0;
		end

reg Pass_300;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_300<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1871==mem[300])&&(Pass_299))
				Pass_300<=1;
			else
				Pass_300<=0;
		end

reg Pass_301;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_301<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1881==mem[301])&&(Pass_300))
				Pass_301<=1;
			else
				Pass_301<=0;
		end

reg Pass_302;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_302<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1891==mem[302])&&(Pass_301))
				Pass_302<=1;
			else
				Pass_302<=0;
		end

reg Pass_303;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_303<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18A1==mem[303])&&(Pass_302))
				Pass_303<=1;
			else
				Pass_303<=0;
		end

reg Pass_304;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_304<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18B1==mem[304])&&(Pass_303))
				Pass_304<=1;
			else
				Pass_304<=0;
		end

reg Pass_305;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_305<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18C1==mem[305])&&(Pass_304))
				Pass_305<=1;
			else
				Pass_305<=0;
		end

reg Pass_306;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_306<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18D1==mem[306])&&(Pass_305))
				Pass_306<=1;
			else
				Pass_306<=0;
		end

reg Pass_307;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_307<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18E1==mem[307])&&(Pass_306))
				Pass_307<=1;
			else
				Pass_307<=0;
		end

reg Pass_308;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_308<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1911==mem[308])&&(Pass_307))
				Pass_308<=1;
			else
				Pass_308<=0;
		end

reg Pass_309;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_309<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1921==mem[309])&&(Pass_308))
				Pass_309<=1;
			else
				Pass_309<=0;
		end

reg Pass_310;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_310<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1931==mem[310])&&(Pass_309))
				Pass_310<=1;
			else
				Pass_310<=0;
		end

reg Pass_311;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_311<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1941==mem[311])&&(Pass_310))
				Pass_311<=1;
			else
				Pass_311<=0;
		end

reg Pass_312;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_312<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1951==mem[312])&&(Pass_311))
				Pass_312<=1;
			else
				Pass_312<=0;
		end

reg Pass_313;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_313<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1961==mem[313])&&(Pass_312))
				Pass_313<=1;
			else
				Pass_313<=0;
		end

reg Pass_314;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_314<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1971==mem[314])&&(Pass_313))
				Pass_314<=1;
			else
				Pass_314<=0;
		end

reg Pass_315;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_315<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1981==mem[315])&&(Pass_314))
				Pass_315<=1;
			else
				Pass_315<=0;
		end

reg Pass_316;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_316<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1991==mem[316])&&(Pass_315))
				Pass_316<=1;
			else
				Pass_316<=0;
		end

reg Pass_317;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_317<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19A1==mem[317])&&(Pass_316))
				Pass_317<=1;
			else
				Pass_317<=0;
		end

reg Pass_318;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_318<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19B1==mem[318])&&(Pass_317))
				Pass_318<=1;
			else
				Pass_318<=0;
		end

reg Pass_319;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_319<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19C1==mem[319])&&(Pass_318))
				Pass_319<=1;
			else
				Pass_319<=0;
		end

reg Pass_320;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_320<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19D1==mem[320])&&(Pass_319))
				Pass_320<=1;
			else
				Pass_320<=0;
		end

reg Pass_321;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_321<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19E1==mem[321])&&(Pass_320))
				Pass_321<=1;
			else
				Pass_321<=0;
		end

reg Pass_322;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_322<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A11==mem[322])&&(Pass_321))
				Pass_322<=1;
			else
				Pass_322<=0;
		end

reg Pass_323;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_323<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A21==mem[323])&&(Pass_322))
				Pass_323<=1;
			else
				Pass_323<=0;
		end

reg Pass_324;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_324<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A31==mem[324])&&(Pass_323))
				Pass_324<=1;
			else
				Pass_324<=0;
		end

reg Pass_325;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_325<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A41==mem[325])&&(Pass_324))
				Pass_325<=1;
			else
				Pass_325<=0;
		end

reg Pass_326;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_326<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A51==mem[326])&&(Pass_325))
				Pass_326<=1;
			else
				Pass_326<=0;
		end

reg Pass_327;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_327<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A61==mem[327])&&(Pass_326))
				Pass_327<=1;
			else
				Pass_327<=0;
		end

reg Pass_328;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_328<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A71==mem[328])&&(Pass_327))
				Pass_328<=1;
			else
				Pass_328<=0;
		end

reg Pass_329;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_329<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A81==mem[329])&&(Pass_328))
				Pass_329<=1;
			else
				Pass_329<=0;
		end

reg Pass_330;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_330<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A91==mem[330])&&(Pass_329))
				Pass_330<=1;
			else
				Pass_330<=0;
		end

reg Pass_331;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_331<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AA1==mem[331])&&(Pass_330))
				Pass_331<=1;
			else
				Pass_331<=0;
		end

reg Pass_332;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_332<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AB1==mem[332])&&(Pass_331))
				Pass_332<=1;
			else
				Pass_332<=0;
		end

reg Pass_333;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_333<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AC1==mem[333])&&(Pass_332))
				Pass_333<=1;
			else
				Pass_333<=0;
		end

reg Pass_334;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_334<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AD1==mem[334])&&(Pass_333))
				Pass_334<=1;
			else
				Pass_334<=0;
		end

reg Pass_335;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_335<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AE1==mem[335])&&(Pass_334))
				Pass_335<=1;
			else
				Pass_335<=0;
		end

reg Pass_336;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_336<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B11==mem[336])&&(Pass_335))
				Pass_336<=1;
			else
				Pass_336<=0;
		end

reg Pass_337;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_337<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B21==mem[337])&&(Pass_336))
				Pass_337<=1;
			else
				Pass_337<=0;
		end

reg Pass_338;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_338<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B31==mem[338])&&(Pass_337))
				Pass_338<=1;
			else
				Pass_338<=0;
		end

reg Pass_339;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_339<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B41==mem[339])&&(Pass_338))
				Pass_339<=1;
			else
				Pass_339<=0;
		end

reg Pass_340;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_340<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B51==mem[340])&&(Pass_339))
				Pass_340<=1;
			else
				Pass_340<=0;
		end

reg Pass_341;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_341<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B61==mem[341])&&(Pass_340))
				Pass_341<=1;
			else
				Pass_341<=0;
		end

reg Pass_342;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_342<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B71==mem[342])&&(Pass_341))
				Pass_342<=1;
			else
				Pass_342<=0;
		end

reg Pass_343;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_343<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B81==mem[343])&&(Pass_342))
				Pass_343<=1;
			else
				Pass_343<=0;
		end

reg Pass_344;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_344<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B91==mem[344])&&(Pass_343))
				Pass_344<=1;
			else
				Pass_344<=0;
		end

reg Pass_345;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_345<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BA1==mem[345])&&(Pass_344))
				Pass_345<=1;
			else
				Pass_345<=0;
		end

reg Pass_346;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_346<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BB1==mem[346])&&(Pass_345))
				Pass_346<=1;
			else
				Pass_346<=0;
		end

reg Pass_347;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_347<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BC1==mem[347])&&(Pass_346))
				Pass_347<=1;
			else
				Pass_347<=0;
		end

reg Pass_348;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_348<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BD1==mem[348])&&(Pass_347))
				Pass_348<=1;
			else
				Pass_348<=0;
		end

reg Pass_349;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_349<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BE1==mem[349])&&(Pass_348))
				Pass_349<=1;
			else
				Pass_349<=0;
		end

reg Pass_350;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_350<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C11==mem[350])&&(Pass_349))
				Pass_350<=1;
			else
				Pass_350<=0;
		end

reg Pass_351;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_351<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C21==mem[351])&&(Pass_350))
				Pass_351<=1;
			else
				Pass_351<=0;
		end

reg Pass_352;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_352<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C31==mem[352])&&(Pass_351))
				Pass_352<=1;
			else
				Pass_352<=0;
		end

reg Pass_353;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_353<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C41==mem[353])&&(Pass_352))
				Pass_353<=1;
			else
				Pass_353<=0;
		end

reg Pass_354;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_354<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C51==mem[354])&&(Pass_353))
				Pass_354<=1;
			else
				Pass_354<=0;
		end

reg Pass_355;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_355<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C61==mem[355])&&(Pass_354))
				Pass_355<=1;
			else
				Pass_355<=0;
		end

reg Pass_356;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_356<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C71==mem[356])&&(Pass_355))
				Pass_356<=1;
			else
				Pass_356<=0;
		end

reg Pass_357;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_357<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C81==mem[357])&&(Pass_356))
				Pass_357<=1;
			else
				Pass_357<=0;
		end

reg Pass_358;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_358<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C91==mem[358])&&(Pass_357))
				Pass_358<=1;
			else
				Pass_358<=0;
		end

reg Pass_359;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_359<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CA1==mem[359])&&(Pass_358))
				Pass_359<=1;
			else
				Pass_359<=0;
		end

reg Pass_360;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_360<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CB1==mem[360])&&(Pass_359))
				Pass_360<=1;
			else
				Pass_360<=0;
		end

reg Pass_361;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_361<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CC1==mem[361])&&(Pass_360))
				Pass_361<=1;
			else
				Pass_361<=0;
		end

reg Pass_362;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_362<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CD1==mem[362])&&(Pass_361))
				Pass_362<=1;
			else
				Pass_362<=0;
		end

reg Pass_363;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_363<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CE1==mem[363])&&(Pass_362))
				Pass_363<=1;
			else
				Pass_363<=0;
		end

reg Pass_364;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_364<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D11==mem[364])&&(Pass_363))
				Pass_364<=1;
			else
				Pass_364<=0;
		end

reg Pass_365;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_365<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D21==mem[365])&&(Pass_364))
				Pass_365<=1;
			else
				Pass_365<=0;
		end

reg Pass_366;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_366<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D31==mem[366])&&(Pass_365))
				Pass_366<=1;
			else
				Pass_366<=0;
		end

reg Pass_367;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_367<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D41==mem[367])&&(Pass_366))
				Pass_367<=1;
			else
				Pass_367<=0;
		end

reg Pass_368;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_368<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D51==mem[368])&&(Pass_367))
				Pass_368<=1;
			else
				Pass_368<=0;
		end

reg Pass_369;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_369<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D61==mem[369])&&(Pass_368))
				Pass_369<=1;
			else
				Pass_369<=0;
		end

reg Pass_370;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_370<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D71==mem[370])&&(Pass_369))
				Pass_370<=1;
			else
				Pass_370<=0;
		end

reg Pass_371;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_371<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D81==mem[371])&&(Pass_370))
				Pass_371<=1;
			else
				Pass_371<=0;
		end

reg Pass_372;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_372<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D91==mem[372])&&(Pass_371))
				Pass_372<=1;
			else
				Pass_372<=0;
		end

reg Pass_373;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_373<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DA1==mem[373])&&(Pass_372))
				Pass_373<=1;
			else
				Pass_373<=0;
		end

reg Pass_374;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_374<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DB1==mem[374])&&(Pass_373))
				Pass_374<=1;
			else
				Pass_374<=0;
		end

reg Pass_375;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_375<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DC1==mem[375])&&(Pass_374))
				Pass_375<=1;
			else
				Pass_375<=0;
		end

reg Pass_376;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_376<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DD1==mem[376])&&(Pass_375))
				Pass_376<=1;
			else
				Pass_376<=0;
		end

reg Pass_377;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_377<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DE1==mem[377])&&(Pass_376))
				Pass_377<=1;
			else
				Pass_377<=0;
		end

reg Pass_378;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_378<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E11==mem[378])&&(Pass_377))
				Pass_378<=1;
			else
				Pass_378<=0;
		end

reg Pass_379;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_379<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E21==mem[379])&&(Pass_378))
				Pass_379<=1;
			else
				Pass_379<=0;
		end

reg Pass_380;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_380<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E31==mem[380])&&(Pass_379))
				Pass_380<=1;
			else
				Pass_380<=0;
		end

reg Pass_381;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_381<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E41==mem[381])&&(Pass_380))
				Pass_381<=1;
			else
				Pass_381<=0;
		end

reg Pass_382;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_382<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E51==mem[382])&&(Pass_381))
				Pass_382<=1;
			else
				Pass_382<=0;
		end

reg Pass_383;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_383<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E61==mem[383])&&(Pass_382))
				Pass_383<=1;
			else
				Pass_383<=0;
		end

reg Pass_384;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_384<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E71==mem[384])&&(Pass_383))
				Pass_384<=1;
			else
				Pass_384<=0;
		end

reg Pass_385;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_385<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E81==mem[385])&&(Pass_384))
				Pass_385<=1;
			else
				Pass_385<=0;
		end

reg Pass_386;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_386<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E91==mem[386])&&(Pass_385))
				Pass_386<=1;
			else
				Pass_386<=0;
		end

reg Pass_387;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_387<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1EA1==mem[387])&&(Pass_386))
				Pass_387<=1;
			else
				Pass_387<=0;
		end

reg Pass_388;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_388<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1EB1==mem[388])&&(Pass_387))
				Pass_388<=1;
			else
				Pass_388<=0;
		end

reg Pass_389;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_389<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1EC1==mem[389])&&(Pass_388))
				Pass_389<=1;
			else
				Pass_389<=0;
		end

reg Pass_390;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_390<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1ED1==mem[390])&&(Pass_389))
				Pass_390<=1;
			else
				Pass_390<=0;
		end

reg Pass_391;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_391<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1EE1==mem[391])&&(Pass_390))
				Pass_391<=1;
			else
				Pass_391<=0;
		end

reg Pass_392;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_392<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1112==mem[392])&&(Pass_391))
				Pass_392<=1;
			else
				Pass_392<=0;
		end

reg Pass_393;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_393<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1122==mem[393])&&(Pass_392))
				Pass_393<=1;
			else
				Pass_393<=0;
		end

reg Pass_394;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_394<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1132==mem[394])&&(Pass_393))
				Pass_394<=1;
			else
				Pass_394<=0;
		end

reg Pass_395;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_395<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1142==mem[395])&&(Pass_394))
				Pass_395<=1;
			else
				Pass_395<=0;
		end

reg Pass_396;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_396<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1152==mem[396])&&(Pass_395))
				Pass_396<=1;
			else
				Pass_396<=0;
		end

reg Pass_397;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_397<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1162==mem[397])&&(Pass_396))
				Pass_397<=1;
			else
				Pass_397<=0;
		end

reg Pass_398;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_398<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1172==mem[398])&&(Pass_397))
				Pass_398<=1;
			else
				Pass_398<=0;
		end

reg Pass_399;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_399<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1182==mem[399])&&(Pass_398))
				Pass_399<=1;
			else
				Pass_399<=0;
		end

reg Pass_400;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_400<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1192==mem[400])&&(Pass_399))
				Pass_400<=1;
			else
				Pass_400<=0;
		end

reg Pass_401;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_401<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11A2==mem[401])&&(Pass_400))
				Pass_401<=1;
			else
				Pass_401<=0;
		end

reg Pass_402;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_402<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11B2==mem[402])&&(Pass_401))
				Pass_402<=1;
			else
				Pass_402<=0;
		end

reg Pass_403;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_403<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11C2==mem[403])&&(Pass_402))
				Pass_403<=1;
			else
				Pass_403<=0;
		end

reg Pass_404;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_404<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11D2==mem[404])&&(Pass_403))
				Pass_404<=1;
			else
				Pass_404<=0;
		end

reg Pass_405;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_405<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11E2==mem[405])&&(Pass_404))
				Pass_405<=1;
			else
				Pass_405<=0;
		end

reg Pass_406;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_406<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1212==mem[406])&&(Pass_405))
				Pass_406<=1;
			else
				Pass_406<=0;
		end

reg Pass_407;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_407<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1222==mem[407])&&(Pass_406))
				Pass_407<=1;
			else
				Pass_407<=0;
		end

reg Pass_408;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_408<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1232==mem[408])&&(Pass_407))
				Pass_408<=1;
			else
				Pass_408<=0;
		end

reg Pass_409;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_409<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1242==mem[409])&&(Pass_408))
				Pass_409<=1;
			else
				Pass_409<=0;
		end

reg Pass_410;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_410<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1252==mem[410])&&(Pass_409))
				Pass_410<=1;
			else
				Pass_410<=0;
		end

reg Pass_411;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_411<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1262==mem[411])&&(Pass_410))
				Pass_411<=1;
			else
				Pass_411<=0;
		end

reg Pass_412;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_412<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1272==mem[412])&&(Pass_411))
				Pass_412<=1;
			else
				Pass_412<=0;
		end

reg Pass_413;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_413<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1282==mem[413])&&(Pass_412))
				Pass_413<=1;
			else
				Pass_413<=0;
		end

reg Pass_414;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_414<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1292==mem[414])&&(Pass_413))
				Pass_414<=1;
			else
				Pass_414<=0;
		end

reg Pass_415;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_415<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12A2==mem[415])&&(Pass_414))
				Pass_415<=1;
			else
				Pass_415<=0;
		end

reg Pass_416;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_416<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12B2==mem[416])&&(Pass_415))
				Pass_416<=1;
			else
				Pass_416<=0;
		end

reg Pass_417;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_417<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12C2==mem[417])&&(Pass_416))
				Pass_417<=1;
			else
				Pass_417<=0;
		end

reg Pass_418;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_418<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12D2==mem[418])&&(Pass_417))
				Pass_418<=1;
			else
				Pass_418<=0;
		end

reg Pass_419;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_419<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12E2==mem[419])&&(Pass_418))
				Pass_419<=1;
			else
				Pass_419<=0;
		end

reg Pass_420;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_420<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1312==mem[420])&&(Pass_419))
				Pass_420<=1;
			else
				Pass_420<=0;
		end

reg Pass_421;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_421<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1322==mem[421])&&(Pass_420))
				Pass_421<=1;
			else
				Pass_421<=0;
		end

reg Pass_422;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_422<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1332==mem[422])&&(Pass_421))
				Pass_422<=1;
			else
				Pass_422<=0;
		end

reg Pass_423;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_423<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1342==mem[423])&&(Pass_422))
				Pass_423<=1;
			else
				Pass_423<=0;
		end

reg Pass_424;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_424<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1352==mem[424])&&(Pass_423))
				Pass_424<=1;
			else
				Pass_424<=0;
		end

reg Pass_425;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_425<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1362==mem[425])&&(Pass_424))
				Pass_425<=1;
			else
				Pass_425<=0;
		end

reg Pass_426;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_426<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1372==mem[426])&&(Pass_425))
				Pass_426<=1;
			else
				Pass_426<=0;
		end

reg Pass_427;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_427<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1382==mem[427])&&(Pass_426))
				Pass_427<=1;
			else
				Pass_427<=0;
		end

reg Pass_428;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_428<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1392==mem[428])&&(Pass_427))
				Pass_428<=1;
			else
				Pass_428<=0;
		end

reg Pass_429;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_429<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13A2==mem[429])&&(Pass_428))
				Pass_429<=1;
			else
				Pass_429<=0;
		end

reg Pass_430;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_430<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13B2==mem[430])&&(Pass_429))
				Pass_430<=1;
			else
				Pass_430<=0;
		end

reg Pass_431;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_431<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13C2==mem[431])&&(Pass_430))
				Pass_431<=1;
			else
				Pass_431<=0;
		end

reg Pass_432;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_432<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13D2==mem[432])&&(Pass_431))
				Pass_432<=1;
			else
				Pass_432<=0;
		end

reg Pass_433;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_433<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13E2==mem[433])&&(Pass_432))
				Pass_433<=1;
			else
				Pass_433<=0;
		end

reg Pass_434;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_434<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1412==mem[434])&&(Pass_433))
				Pass_434<=1;
			else
				Pass_434<=0;
		end

reg Pass_435;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_435<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1422==mem[435])&&(Pass_434))
				Pass_435<=1;
			else
				Pass_435<=0;
		end

reg Pass_436;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_436<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1432==mem[436])&&(Pass_435))
				Pass_436<=1;
			else
				Pass_436<=0;
		end

reg Pass_437;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_437<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1442==mem[437])&&(Pass_436))
				Pass_437<=1;
			else
				Pass_437<=0;
		end

reg Pass_438;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_438<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1452==mem[438])&&(Pass_437))
				Pass_438<=1;
			else
				Pass_438<=0;
		end

reg Pass_439;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_439<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1462==mem[439])&&(Pass_438))
				Pass_439<=1;
			else
				Pass_439<=0;
		end

reg Pass_440;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_440<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1472==mem[440])&&(Pass_439))
				Pass_440<=1;
			else
				Pass_440<=0;
		end

reg Pass_441;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_441<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1482==mem[441])&&(Pass_440))
				Pass_441<=1;
			else
				Pass_441<=0;
		end

reg Pass_442;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_442<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1492==mem[442])&&(Pass_441))
				Pass_442<=1;
			else
				Pass_442<=0;
		end

reg Pass_443;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_443<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14A2==mem[443])&&(Pass_442))
				Pass_443<=1;
			else
				Pass_443<=0;
		end

reg Pass_444;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_444<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14B2==mem[444])&&(Pass_443))
				Pass_444<=1;
			else
				Pass_444<=0;
		end

reg Pass_445;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_445<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14C2==mem[445])&&(Pass_444))
				Pass_445<=1;
			else
				Pass_445<=0;
		end

reg Pass_446;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_446<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14D2==mem[446])&&(Pass_445))
				Pass_446<=1;
			else
				Pass_446<=0;
		end

reg Pass_447;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_447<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14E2==mem[447])&&(Pass_446))
				Pass_447<=1;
			else
				Pass_447<=0;
		end

reg Pass_448;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_448<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1512==mem[448])&&(Pass_447))
				Pass_448<=1;
			else
				Pass_448<=0;
		end

reg Pass_449;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_449<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1522==mem[449])&&(Pass_448))
				Pass_449<=1;
			else
				Pass_449<=0;
		end

reg Pass_450;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_450<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1532==mem[450])&&(Pass_449))
				Pass_450<=1;
			else
				Pass_450<=0;
		end

reg Pass_451;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_451<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1542==mem[451])&&(Pass_450))
				Pass_451<=1;
			else
				Pass_451<=0;
		end

reg Pass_452;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_452<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1552==mem[452])&&(Pass_451))
				Pass_452<=1;
			else
				Pass_452<=0;
		end

reg Pass_453;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_453<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1562==mem[453])&&(Pass_452))
				Pass_453<=1;
			else
				Pass_453<=0;
		end

reg Pass_454;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_454<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1572==mem[454])&&(Pass_453))
				Pass_454<=1;
			else
				Pass_454<=0;
		end

reg Pass_455;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_455<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1582==mem[455])&&(Pass_454))
				Pass_455<=1;
			else
				Pass_455<=0;
		end

reg Pass_456;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_456<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1592==mem[456])&&(Pass_455))
				Pass_456<=1;
			else
				Pass_456<=0;
		end

reg Pass_457;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_457<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15A2==mem[457])&&(Pass_456))
				Pass_457<=1;
			else
				Pass_457<=0;
		end

reg Pass_458;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_458<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15B2==mem[458])&&(Pass_457))
				Pass_458<=1;
			else
				Pass_458<=0;
		end

reg Pass_459;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_459<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15C2==mem[459])&&(Pass_458))
				Pass_459<=1;
			else
				Pass_459<=0;
		end

reg Pass_460;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_460<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15D2==mem[460])&&(Pass_459))
				Pass_460<=1;
			else
				Pass_460<=0;
		end

reg Pass_461;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_461<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15E2==mem[461])&&(Pass_460))
				Pass_461<=1;
			else
				Pass_461<=0;
		end

reg Pass_462;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_462<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1612==mem[462])&&(Pass_461))
				Pass_462<=1;
			else
				Pass_462<=0;
		end

reg Pass_463;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_463<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1622==mem[463])&&(Pass_462))
				Pass_463<=1;
			else
				Pass_463<=0;
		end

reg Pass_464;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_464<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1632==mem[464])&&(Pass_463))
				Pass_464<=1;
			else
				Pass_464<=0;
		end

reg Pass_465;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_465<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1642==mem[465])&&(Pass_464))
				Pass_465<=1;
			else
				Pass_465<=0;
		end

reg Pass_466;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_466<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1652==mem[466])&&(Pass_465))
				Pass_466<=1;
			else
				Pass_466<=0;
		end

reg Pass_467;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_467<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1662==mem[467])&&(Pass_466))
				Pass_467<=1;
			else
				Pass_467<=0;
		end

reg Pass_468;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_468<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1672==mem[468])&&(Pass_467))
				Pass_468<=1;
			else
				Pass_468<=0;
		end

reg Pass_469;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_469<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1682==mem[469])&&(Pass_468))
				Pass_469<=1;
			else
				Pass_469<=0;
		end

reg Pass_470;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_470<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1692==mem[470])&&(Pass_469))
				Pass_470<=1;
			else
				Pass_470<=0;
		end

reg Pass_471;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_471<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16A2==mem[471])&&(Pass_470))
				Pass_471<=1;
			else
				Pass_471<=0;
		end

reg Pass_472;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_472<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16B2==mem[472])&&(Pass_471))
				Pass_472<=1;
			else
				Pass_472<=0;
		end

reg Pass_473;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_473<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16C2==mem[473])&&(Pass_472))
				Pass_473<=1;
			else
				Pass_473<=0;
		end

reg Pass_474;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_474<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16D2==mem[474])&&(Pass_473))
				Pass_474<=1;
			else
				Pass_474<=0;
		end

reg Pass_475;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_475<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16E2==mem[475])&&(Pass_474))
				Pass_475<=1;
			else
				Pass_475<=0;
		end

reg Pass_476;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_476<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1712==mem[476])&&(Pass_475))
				Pass_476<=1;
			else
				Pass_476<=0;
		end

reg Pass_477;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_477<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1722==mem[477])&&(Pass_476))
				Pass_477<=1;
			else
				Pass_477<=0;
		end

reg Pass_478;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_478<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1732==mem[478])&&(Pass_477))
				Pass_478<=1;
			else
				Pass_478<=0;
		end

reg Pass_479;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_479<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1742==mem[479])&&(Pass_478))
				Pass_479<=1;
			else
				Pass_479<=0;
		end

reg Pass_480;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_480<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1752==mem[480])&&(Pass_479))
				Pass_480<=1;
			else
				Pass_480<=0;
		end

reg Pass_481;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_481<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1762==mem[481])&&(Pass_480))
				Pass_481<=1;
			else
				Pass_481<=0;
		end

reg Pass_482;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_482<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1772==mem[482])&&(Pass_481))
				Pass_482<=1;
			else
				Pass_482<=0;
		end

reg Pass_483;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_483<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1782==mem[483])&&(Pass_482))
				Pass_483<=1;
			else
				Pass_483<=0;
		end

reg Pass_484;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_484<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1792==mem[484])&&(Pass_483))
				Pass_484<=1;
			else
				Pass_484<=0;
		end

reg Pass_485;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_485<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17A2==mem[485])&&(Pass_484))
				Pass_485<=1;
			else
				Pass_485<=0;
		end

reg Pass_486;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_486<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17B2==mem[486])&&(Pass_485))
				Pass_486<=1;
			else
				Pass_486<=0;
		end

reg Pass_487;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_487<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17C2==mem[487])&&(Pass_486))
				Pass_487<=1;
			else
				Pass_487<=0;
		end

reg Pass_488;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_488<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17D2==mem[488])&&(Pass_487))
				Pass_488<=1;
			else
				Pass_488<=0;
		end

reg Pass_489;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_489<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17E2==mem[489])&&(Pass_488))
				Pass_489<=1;
			else
				Pass_489<=0;
		end

reg Pass_490;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_490<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1812==mem[490])&&(Pass_489))
				Pass_490<=1;
			else
				Pass_490<=0;
		end

reg Pass_491;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_491<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1822==mem[491])&&(Pass_490))
				Pass_491<=1;
			else
				Pass_491<=0;
		end

reg Pass_492;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_492<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1832==mem[492])&&(Pass_491))
				Pass_492<=1;
			else
				Pass_492<=0;
		end

reg Pass_493;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_493<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1842==mem[493])&&(Pass_492))
				Pass_493<=1;
			else
				Pass_493<=0;
		end

reg Pass_494;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_494<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1852==mem[494])&&(Pass_493))
				Pass_494<=1;
			else
				Pass_494<=0;
		end

reg Pass_495;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_495<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1862==mem[495])&&(Pass_494))
				Pass_495<=1;
			else
				Pass_495<=0;
		end

reg Pass_496;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_496<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1872==mem[496])&&(Pass_495))
				Pass_496<=1;
			else
				Pass_496<=0;
		end

reg Pass_497;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_497<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1882==mem[497])&&(Pass_496))
				Pass_497<=1;
			else
				Pass_497<=0;
		end

reg Pass_498;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_498<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1892==mem[498])&&(Pass_497))
				Pass_498<=1;
			else
				Pass_498<=0;
		end

reg Pass_499;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_499<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18A2==mem[499])&&(Pass_498))
				Pass_499<=1;
			else
				Pass_499<=0;
		end

reg Pass_500;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_500<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18B2==mem[500])&&(Pass_499))
				Pass_500<=1;
			else
				Pass_500<=0;
		end

reg Pass_501;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_501<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18C2==mem[501])&&(Pass_500))
				Pass_501<=1;
			else
				Pass_501<=0;
		end

reg Pass_502;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_502<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18D2==mem[502])&&(Pass_501))
				Pass_502<=1;
			else
				Pass_502<=0;
		end

reg Pass_503;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_503<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18E2==mem[503])&&(Pass_502))
				Pass_503<=1;
			else
				Pass_503<=0;
		end

reg Pass_504;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_504<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1912==mem[504])&&(Pass_503))
				Pass_504<=1;
			else
				Pass_504<=0;
		end

reg Pass_505;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_505<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1922==mem[505])&&(Pass_504))
				Pass_505<=1;
			else
				Pass_505<=0;
		end

reg Pass_506;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_506<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1932==mem[506])&&(Pass_505))
				Pass_506<=1;
			else
				Pass_506<=0;
		end

reg Pass_507;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_507<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1942==mem[507])&&(Pass_506))
				Pass_507<=1;
			else
				Pass_507<=0;
		end

reg Pass_508;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_508<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1952==mem[508])&&(Pass_507))
				Pass_508<=1;
			else
				Pass_508<=0;
		end

reg Pass_509;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_509<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1962==mem[509])&&(Pass_508))
				Pass_509<=1;
			else
				Pass_509<=0;
		end

reg Pass_510;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_510<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1972==mem[510])&&(Pass_509))
				Pass_510<=1;
			else
				Pass_510<=0;
		end

reg Pass_511;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_511<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1982==mem[511])&&(Pass_510))
				Pass_511<=1;
			else
				Pass_511<=0;
		end

reg Pass_512;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_512<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1992==mem[512])&&(Pass_511))
				Pass_512<=1;
			else
				Pass_512<=0;
		end

reg Pass_513;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_513<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19A2==mem[513])&&(Pass_512))
				Pass_513<=1;
			else
				Pass_513<=0;
		end

reg Pass_514;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_514<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19B2==mem[514])&&(Pass_513))
				Pass_514<=1;
			else
				Pass_514<=0;
		end

reg Pass_515;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_515<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19C2==mem[515])&&(Pass_514))
				Pass_515<=1;
			else
				Pass_515<=0;
		end

reg Pass_516;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_516<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19D2==mem[516])&&(Pass_515))
				Pass_516<=1;
			else
				Pass_516<=0;
		end

reg Pass_517;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_517<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19E2==mem[517])&&(Pass_516))
				Pass_517<=1;
			else
				Pass_517<=0;
		end

reg Pass_518;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_518<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A12==mem[518])&&(Pass_517))
				Pass_518<=1;
			else
				Pass_518<=0;
		end

reg Pass_519;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_519<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A22==mem[519])&&(Pass_518))
				Pass_519<=1;
			else
				Pass_519<=0;
		end

reg Pass_520;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_520<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A32==mem[520])&&(Pass_519))
				Pass_520<=1;
			else
				Pass_520<=0;
		end

reg Pass_521;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_521<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A42==mem[521])&&(Pass_520))
				Pass_521<=1;
			else
				Pass_521<=0;
		end

reg Pass_522;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_522<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A52==mem[522])&&(Pass_521))
				Pass_522<=1;
			else
				Pass_522<=0;
		end

reg Pass_523;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_523<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A62==mem[523])&&(Pass_522))
				Pass_523<=1;
			else
				Pass_523<=0;
		end

reg Pass_524;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_524<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A72==mem[524])&&(Pass_523))
				Pass_524<=1;
			else
				Pass_524<=0;
		end

reg Pass_525;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_525<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A82==mem[525])&&(Pass_524))
				Pass_525<=1;
			else
				Pass_525<=0;
		end

reg Pass_526;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_526<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A92==mem[526])&&(Pass_525))
				Pass_526<=1;
			else
				Pass_526<=0;
		end

reg Pass_527;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_527<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AA2==mem[527])&&(Pass_526))
				Pass_527<=1;
			else
				Pass_527<=0;
		end

reg Pass_528;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_528<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AB2==mem[528])&&(Pass_527))
				Pass_528<=1;
			else
				Pass_528<=0;
		end

reg Pass_529;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_529<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AC2==mem[529])&&(Pass_528))
				Pass_529<=1;
			else
				Pass_529<=0;
		end

reg Pass_530;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_530<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AD2==mem[530])&&(Pass_529))
				Pass_530<=1;
			else
				Pass_530<=0;
		end

reg Pass_531;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_531<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AE2==mem[531])&&(Pass_530))
				Pass_531<=1;
			else
				Pass_531<=0;
		end

reg Pass_532;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_532<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B12==mem[532])&&(Pass_531))
				Pass_532<=1;
			else
				Pass_532<=0;
		end

reg Pass_533;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_533<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B22==mem[533])&&(Pass_532))
				Pass_533<=1;
			else
				Pass_533<=0;
		end

reg Pass_534;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_534<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B32==mem[534])&&(Pass_533))
				Pass_534<=1;
			else
				Pass_534<=0;
		end

reg Pass_535;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_535<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B42==mem[535])&&(Pass_534))
				Pass_535<=1;
			else
				Pass_535<=0;
		end

reg Pass_536;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_536<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B52==mem[536])&&(Pass_535))
				Pass_536<=1;
			else
				Pass_536<=0;
		end

reg Pass_537;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_537<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B62==mem[537])&&(Pass_536))
				Pass_537<=1;
			else
				Pass_537<=0;
		end

reg Pass_538;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_538<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B72==mem[538])&&(Pass_537))
				Pass_538<=1;
			else
				Pass_538<=0;
		end

reg Pass_539;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_539<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B82==mem[539])&&(Pass_538))
				Pass_539<=1;
			else
				Pass_539<=0;
		end

reg Pass_540;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_540<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B92==mem[540])&&(Pass_539))
				Pass_540<=1;
			else
				Pass_540<=0;
		end

reg Pass_541;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_541<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BA2==mem[541])&&(Pass_540))
				Pass_541<=1;
			else
				Pass_541<=0;
		end

reg Pass_542;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_542<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BB2==mem[542])&&(Pass_541))
				Pass_542<=1;
			else
				Pass_542<=0;
		end

reg Pass_543;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_543<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BC2==mem[543])&&(Pass_542))
				Pass_543<=1;
			else
				Pass_543<=0;
		end

reg Pass_544;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_544<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BD2==mem[544])&&(Pass_543))
				Pass_544<=1;
			else
				Pass_544<=0;
		end

reg Pass_545;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_545<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BE2==mem[545])&&(Pass_544))
				Pass_545<=1;
			else
				Pass_545<=0;
		end

reg Pass_546;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_546<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C12==mem[546])&&(Pass_545))
				Pass_546<=1;
			else
				Pass_546<=0;
		end

reg Pass_547;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_547<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C22==mem[547])&&(Pass_546))
				Pass_547<=1;
			else
				Pass_547<=0;
		end

reg Pass_548;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_548<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C32==mem[548])&&(Pass_547))
				Pass_548<=1;
			else
				Pass_548<=0;
		end

reg Pass_549;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_549<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C42==mem[549])&&(Pass_548))
				Pass_549<=1;
			else
				Pass_549<=0;
		end

reg Pass_550;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_550<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C52==mem[550])&&(Pass_549))
				Pass_550<=1;
			else
				Pass_550<=0;
		end

reg Pass_551;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_551<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C62==mem[551])&&(Pass_550))
				Pass_551<=1;
			else
				Pass_551<=0;
		end

reg Pass_552;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_552<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C72==mem[552])&&(Pass_551))
				Pass_552<=1;
			else
				Pass_552<=0;
		end

reg Pass_553;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_553<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C82==mem[553])&&(Pass_552))
				Pass_553<=1;
			else
				Pass_553<=0;
		end

reg Pass_554;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_554<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C92==mem[554])&&(Pass_553))
				Pass_554<=1;
			else
				Pass_554<=0;
		end

reg Pass_555;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_555<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CA2==mem[555])&&(Pass_554))
				Pass_555<=1;
			else
				Pass_555<=0;
		end

reg Pass_556;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_556<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CB2==mem[556])&&(Pass_555))
				Pass_556<=1;
			else
				Pass_556<=0;
		end

reg Pass_557;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_557<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CC2==mem[557])&&(Pass_556))
				Pass_557<=1;
			else
				Pass_557<=0;
		end

reg Pass_558;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_558<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CD2==mem[558])&&(Pass_557))
				Pass_558<=1;
			else
				Pass_558<=0;
		end

reg Pass_559;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_559<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CE2==mem[559])&&(Pass_558))
				Pass_559<=1;
			else
				Pass_559<=0;
		end

reg Pass_560;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_560<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D12==mem[560])&&(Pass_559))
				Pass_560<=1;
			else
				Pass_560<=0;
		end

reg Pass_561;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_561<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D22==mem[561])&&(Pass_560))
				Pass_561<=1;
			else
				Pass_561<=0;
		end

reg Pass_562;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_562<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D32==mem[562])&&(Pass_561))
				Pass_562<=1;
			else
				Pass_562<=0;
		end

reg Pass_563;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_563<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D42==mem[563])&&(Pass_562))
				Pass_563<=1;
			else
				Pass_563<=0;
		end

reg Pass_564;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_564<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D52==mem[564])&&(Pass_563))
				Pass_564<=1;
			else
				Pass_564<=0;
		end

reg Pass_565;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_565<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D62==mem[565])&&(Pass_564))
				Pass_565<=1;
			else
				Pass_565<=0;
		end

reg Pass_566;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_566<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D72==mem[566])&&(Pass_565))
				Pass_566<=1;
			else
				Pass_566<=0;
		end

reg Pass_567;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_567<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D82==mem[567])&&(Pass_566))
				Pass_567<=1;
			else
				Pass_567<=0;
		end

reg Pass_568;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_568<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D92==mem[568])&&(Pass_567))
				Pass_568<=1;
			else
				Pass_568<=0;
		end

reg Pass_569;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_569<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DA2==mem[569])&&(Pass_568))
				Pass_569<=1;
			else
				Pass_569<=0;
		end

reg Pass_570;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_570<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DB2==mem[570])&&(Pass_569))
				Pass_570<=1;
			else
				Pass_570<=0;
		end

reg Pass_571;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_571<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DC2==mem[571])&&(Pass_570))
				Pass_571<=1;
			else
				Pass_571<=0;
		end

reg Pass_572;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_572<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DD2==mem[572])&&(Pass_571))
				Pass_572<=1;
			else
				Pass_572<=0;
		end

reg Pass_573;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_573<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DE2==mem[573])&&(Pass_572))
				Pass_573<=1;
			else
				Pass_573<=0;
		end

reg Pass_574;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_574<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E12==mem[574])&&(Pass_573))
				Pass_574<=1;
			else
				Pass_574<=0;
		end

reg Pass_575;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_575<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E22==mem[575])&&(Pass_574))
				Pass_575<=1;
			else
				Pass_575<=0;
		end

reg Pass_576;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_576<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E32==mem[576])&&(Pass_575))
				Pass_576<=1;
			else
				Pass_576<=0;
		end

reg Pass_577;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_577<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E42==mem[577])&&(Pass_576))
				Pass_577<=1;
			else
				Pass_577<=0;
		end

reg Pass_578;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_578<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E52==mem[578])&&(Pass_577))
				Pass_578<=1;
			else
				Pass_578<=0;
		end

reg Pass_579;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_579<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E62==mem[579])&&(Pass_578))
				Pass_579<=1;
			else
				Pass_579<=0;
		end

reg Pass_580;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_580<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E72==mem[580])&&(Pass_579))
				Pass_580<=1;
			else
				Pass_580<=0;
		end

reg Pass_581;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_581<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E82==mem[581])&&(Pass_580))
				Pass_581<=1;
			else
				Pass_581<=0;
		end

reg Pass_582;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_582<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E92==mem[582])&&(Pass_581))
				Pass_582<=1;
			else
				Pass_582<=0;
		end

reg Pass_583;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_583<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1EA2==mem[583])&&(Pass_582))
				Pass_583<=1;
			else
				Pass_583<=0;
		end

reg Pass_584;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_584<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1EB2==mem[584])&&(Pass_583))
				Pass_584<=1;
			else
				Pass_584<=0;
		end

reg Pass_585;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_585<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1EC2==mem[585])&&(Pass_584))
				Pass_585<=1;
			else
				Pass_585<=0;
		end

reg Pass_586;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_586<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1ED2==mem[586])&&(Pass_585))
				Pass_586<=1;
			else
				Pass_586<=0;
		end

reg Pass_587;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_587<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1EE2==mem[587])&&(Pass_586))
				Pass_587<=1;
			else
				Pass_587<=0;
		end

reg Pass_588;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_588<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1113==mem[588])&&(Pass_587))
				Pass_588<=1;
			else
				Pass_588<=0;
		end

reg Pass_589;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_589<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1123==mem[589])&&(Pass_588))
				Pass_589<=1;
			else
				Pass_589<=0;
		end

reg Pass_590;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_590<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1133==mem[590])&&(Pass_589))
				Pass_590<=1;
			else
				Pass_590<=0;
		end

reg Pass_591;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_591<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1143==mem[591])&&(Pass_590))
				Pass_591<=1;
			else
				Pass_591<=0;
		end

reg Pass_592;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_592<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1153==mem[592])&&(Pass_591))
				Pass_592<=1;
			else
				Pass_592<=0;
		end

reg Pass_593;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_593<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1163==mem[593])&&(Pass_592))
				Pass_593<=1;
			else
				Pass_593<=0;
		end

reg Pass_594;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_594<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1173==mem[594])&&(Pass_593))
				Pass_594<=1;
			else
				Pass_594<=0;
		end

reg Pass_595;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_595<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1183==mem[595])&&(Pass_594))
				Pass_595<=1;
			else
				Pass_595<=0;
		end

reg Pass_596;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_596<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1193==mem[596])&&(Pass_595))
				Pass_596<=1;
			else
				Pass_596<=0;
		end

reg Pass_597;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_597<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11A3==mem[597])&&(Pass_596))
				Pass_597<=1;
			else
				Pass_597<=0;
		end

reg Pass_598;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_598<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11B3==mem[598])&&(Pass_597))
				Pass_598<=1;
			else
				Pass_598<=0;
		end

reg Pass_599;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_599<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11C3==mem[599])&&(Pass_598))
				Pass_599<=1;
			else
				Pass_599<=0;
		end

reg Pass_600;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_600<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11D3==mem[600])&&(Pass_599))
				Pass_600<=1;
			else
				Pass_600<=0;
		end

reg Pass_601;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_601<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P11E3==mem[601])&&(Pass_600))
				Pass_601<=1;
			else
				Pass_601<=0;
		end

reg Pass_602;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_602<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1213==mem[602])&&(Pass_601))
				Pass_602<=1;
			else
				Pass_602<=0;
		end

reg Pass_603;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_603<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1223==mem[603])&&(Pass_602))
				Pass_603<=1;
			else
				Pass_603<=0;
		end

reg Pass_604;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_604<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1233==mem[604])&&(Pass_603))
				Pass_604<=1;
			else
				Pass_604<=0;
		end

reg Pass_605;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_605<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1243==mem[605])&&(Pass_604))
				Pass_605<=1;
			else
				Pass_605<=0;
		end

reg Pass_606;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_606<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1253==mem[606])&&(Pass_605))
				Pass_606<=1;
			else
				Pass_606<=0;
		end

reg Pass_607;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_607<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1263==mem[607])&&(Pass_606))
				Pass_607<=1;
			else
				Pass_607<=0;
		end

reg Pass_608;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_608<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1273==mem[608])&&(Pass_607))
				Pass_608<=1;
			else
				Pass_608<=0;
		end

reg Pass_609;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_609<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1283==mem[609])&&(Pass_608))
				Pass_609<=1;
			else
				Pass_609<=0;
		end

reg Pass_610;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_610<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1293==mem[610])&&(Pass_609))
				Pass_610<=1;
			else
				Pass_610<=0;
		end

reg Pass_611;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_611<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12A3==mem[611])&&(Pass_610))
				Pass_611<=1;
			else
				Pass_611<=0;
		end

reg Pass_612;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_612<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12B3==mem[612])&&(Pass_611))
				Pass_612<=1;
			else
				Pass_612<=0;
		end

reg Pass_613;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_613<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12C3==mem[613])&&(Pass_612))
				Pass_613<=1;
			else
				Pass_613<=0;
		end

reg Pass_614;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_614<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12D3==mem[614])&&(Pass_613))
				Pass_614<=1;
			else
				Pass_614<=0;
		end

reg Pass_615;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_615<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P12E3==mem[615])&&(Pass_614))
				Pass_615<=1;
			else
				Pass_615<=0;
		end

reg Pass_616;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_616<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1313==mem[616])&&(Pass_615))
				Pass_616<=1;
			else
				Pass_616<=0;
		end

reg Pass_617;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_617<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1323==mem[617])&&(Pass_616))
				Pass_617<=1;
			else
				Pass_617<=0;
		end

reg Pass_618;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_618<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1333==mem[618])&&(Pass_617))
				Pass_618<=1;
			else
				Pass_618<=0;
		end

reg Pass_619;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_619<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1343==mem[619])&&(Pass_618))
				Pass_619<=1;
			else
				Pass_619<=0;
		end

reg Pass_620;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_620<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1353==mem[620])&&(Pass_619))
				Pass_620<=1;
			else
				Pass_620<=0;
		end

reg Pass_621;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_621<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1363==mem[621])&&(Pass_620))
				Pass_621<=1;
			else
				Pass_621<=0;
		end

reg Pass_622;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_622<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1373==mem[622])&&(Pass_621))
				Pass_622<=1;
			else
				Pass_622<=0;
		end

reg Pass_623;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_623<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1383==mem[623])&&(Pass_622))
				Pass_623<=1;
			else
				Pass_623<=0;
		end

reg Pass_624;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_624<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1393==mem[624])&&(Pass_623))
				Pass_624<=1;
			else
				Pass_624<=0;
		end

reg Pass_625;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_625<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13A3==mem[625])&&(Pass_624))
				Pass_625<=1;
			else
				Pass_625<=0;
		end

reg Pass_626;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_626<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13B3==mem[626])&&(Pass_625))
				Pass_626<=1;
			else
				Pass_626<=0;
		end

reg Pass_627;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_627<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13C3==mem[627])&&(Pass_626))
				Pass_627<=1;
			else
				Pass_627<=0;
		end

reg Pass_628;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_628<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13D3==mem[628])&&(Pass_627))
				Pass_628<=1;
			else
				Pass_628<=0;
		end

reg Pass_629;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_629<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P13E3==mem[629])&&(Pass_628))
				Pass_629<=1;
			else
				Pass_629<=0;
		end

reg Pass_630;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_630<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1413==mem[630])&&(Pass_629))
				Pass_630<=1;
			else
				Pass_630<=0;
		end

reg Pass_631;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_631<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1423==mem[631])&&(Pass_630))
				Pass_631<=1;
			else
				Pass_631<=0;
		end

reg Pass_632;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_632<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1433==mem[632])&&(Pass_631))
				Pass_632<=1;
			else
				Pass_632<=0;
		end

reg Pass_633;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_633<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1443==mem[633])&&(Pass_632))
				Pass_633<=1;
			else
				Pass_633<=0;
		end

reg Pass_634;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_634<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1453==mem[634])&&(Pass_633))
				Pass_634<=1;
			else
				Pass_634<=0;
		end

reg Pass_635;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_635<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1463==mem[635])&&(Pass_634))
				Pass_635<=1;
			else
				Pass_635<=0;
		end

reg Pass_636;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_636<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1473==mem[636])&&(Pass_635))
				Pass_636<=1;
			else
				Pass_636<=0;
		end

reg Pass_637;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_637<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1483==mem[637])&&(Pass_636))
				Pass_637<=1;
			else
				Pass_637<=0;
		end

reg Pass_638;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_638<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1493==mem[638])&&(Pass_637))
				Pass_638<=1;
			else
				Pass_638<=0;
		end

reg Pass_639;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_639<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14A3==mem[639])&&(Pass_638))
				Pass_639<=1;
			else
				Pass_639<=0;
		end

reg Pass_640;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_640<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14B3==mem[640])&&(Pass_639))
				Pass_640<=1;
			else
				Pass_640<=0;
		end

reg Pass_641;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_641<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14C3==mem[641])&&(Pass_640))
				Pass_641<=1;
			else
				Pass_641<=0;
		end

reg Pass_642;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_642<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14D3==mem[642])&&(Pass_641))
				Pass_642<=1;
			else
				Pass_642<=0;
		end

reg Pass_643;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_643<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P14E3==mem[643])&&(Pass_642))
				Pass_643<=1;
			else
				Pass_643<=0;
		end

reg Pass_644;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_644<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1513==mem[644])&&(Pass_643))
				Pass_644<=1;
			else
				Pass_644<=0;
		end

reg Pass_645;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_645<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1523==mem[645])&&(Pass_644))
				Pass_645<=1;
			else
				Pass_645<=0;
		end

reg Pass_646;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_646<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1533==mem[646])&&(Pass_645))
				Pass_646<=1;
			else
				Pass_646<=0;
		end

reg Pass_647;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_647<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1543==mem[647])&&(Pass_646))
				Pass_647<=1;
			else
				Pass_647<=0;
		end

reg Pass_648;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_648<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1553==mem[648])&&(Pass_647))
				Pass_648<=1;
			else
				Pass_648<=0;
		end

reg Pass_649;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_649<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1563==mem[649])&&(Pass_648))
				Pass_649<=1;
			else
				Pass_649<=0;
		end

reg Pass_650;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_650<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1573==mem[650])&&(Pass_649))
				Pass_650<=1;
			else
				Pass_650<=0;
		end

reg Pass_651;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_651<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1583==mem[651])&&(Pass_650))
				Pass_651<=1;
			else
				Pass_651<=0;
		end

reg Pass_652;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_652<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1593==mem[652])&&(Pass_651))
				Pass_652<=1;
			else
				Pass_652<=0;
		end

reg Pass_653;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_653<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15A3==mem[653])&&(Pass_652))
				Pass_653<=1;
			else
				Pass_653<=0;
		end

reg Pass_654;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_654<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15B3==mem[654])&&(Pass_653))
				Pass_654<=1;
			else
				Pass_654<=0;
		end

reg Pass_655;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_655<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15C3==mem[655])&&(Pass_654))
				Pass_655<=1;
			else
				Pass_655<=0;
		end

reg Pass_656;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_656<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15D3==mem[656])&&(Pass_655))
				Pass_656<=1;
			else
				Pass_656<=0;
		end

reg Pass_657;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_657<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P15E3==mem[657])&&(Pass_656))
				Pass_657<=1;
			else
				Pass_657<=0;
		end

reg Pass_658;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_658<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1613==mem[658])&&(Pass_657))
				Pass_658<=1;
			else
				Pass_658<=0;
		end

reg Pass_659;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_659<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1623==mem[659])&&(Pass_658))
				Pass_659<=1;
			else
				Pass_659<=0;
		end

reg Pass_660;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_660<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1633==mem[660])&&(Pass_659))
				Pass_660<=1;
			else
				Pass_660<=0;
		end

reg Pass_661;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_661<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1643==mem[661])&&(Pass_660))
				Pass_661<=1;
			else
				Pass_661<=0;
		end

reg Pass_662;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_662<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1653==mem[662])&&(Pass_661))
				Pass_662<=1;
			else
				Pass_662<=0;
		end

reg Pass_663;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_663<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1663==mem[663])&&(Pass_662))
				Pass_663<=1;
			else
				Pass_663<=0;
		end

reg Pass_664;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_664<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1673==mem[664])&&(Pass_663))
				Pass_664<=1;
			else
				Pass_664<=0;
		end

reg Pass_665;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_665<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1683==mem[665])&&(Pass_664))
				Pass_665<=1;
			else
				Pass_665<=0;
		end

reg Pass_666;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_666<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1693==mem[666])&&(Pass_665))
				Pass_666<=1;
			else
				Pass_666<=0;
		end

reg Pass_667;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_667<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16A3==mem[667])&&(Pass_666))
				Pass_667<=1;
			else
				Pass_667<=0;
		end

reg Pass_668;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_668<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16B3==mem[668])&&(Pass_667))
				Pass_668<=1;
			else
				Pass_668<=0;
		end

reg Pass_669;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_669<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16C3==mem[669])&&(Pass_668))
				Pass_669<=1;
			else
				Pass_669<=0;
		end

reg Pass_670;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_670<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16D3==mem[670])&&(Pass_669))
				Pass_670<=1;
			else
				Pass_670<=0;
		end

reg Pass_671;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_671<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P16E3==mem[671])&&(Pass_670))
				Pass_671<=1;
			else
				Pass_671<=0;
		end

reg Pass_672;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_672<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1713==mem[672])&&(Pass_671))
				Pass_672<=1;
			else
				Pass_672<=0;
		end

reg Pass_673;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_673<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1723==mem[673])&&(Pass_672))
				Pass_673<=1;
			else
				Pass_673<=0;
		end

reg Pass_674;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_674<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1733==mem[674])&&(Pass_673))
				Pass_674<=1;
			else
				Pass_674<=0;
		end

reg Pass_675;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_675<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1743==mem[675])&&(Pass_674))
				Pass_675<=1;
			else
				Pass_675<=0;
		end

reg Pass_676;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_676<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1753==mem[676])&&(Pass_675))
				Pass_676<=1;
			else
				Pass_676<=0;
		end

reg Pass_677;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_677<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1763==mem[677])&&(Pass_676))
				Pass_677<=1;
			else
				Pass_677<=0;
		end

reg Pass_678;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_678<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1773==mem[678])&&(Pass_677))
				Pass_678<=1;
			else
				Pass_678<=0;
		end

reg Pass_679;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_679<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1783==mem[679])&&(Pass_678))
				Pass_679<=1;
			else
				Pass_679<=0;
		end

reg Pass_680;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_680<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1793==mem[680])&&(Pass_679))
				Pass_680<=1;
			else
				Pass_680<=0;
		end

reg Pass_681;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_681<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17A3==mem[681])&&(Pass_680))
				Pass_681<=1;
			else
				Pass_681<=0;
		end

reg Pass_682;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_682<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17B3==mem[682])&&(Pass_681))
				Pass_682<=1;
			else
				Pass_682<=0;
		end

reg Pass_683;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_683<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17C3==mem[683])&&(Pass_682))
				Pass_683<=1;
			else
				Pass_683<=0;
		end

reg Pass_684;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_684<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17D3==mem[684])&&(Pass_683))
				Pass_684<=1;
			else
				Pass_684<=0;
		end

reg Pass_685;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_685<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P17E3==mem[685])&&(Pass_684))
				Pass_685<=1;
			else
				Pass_685<=0;
		end

reg Pass_686;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_686<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1813==mem[686])&&(Pass_685))
				Pass_686<=1;
			else
				Pass_686<=0;
		end

reg Pass_687;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_687<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1823==mem[687])&&(Pass_686))
				Pass_687<=1;
			else
				Pass_687<=0;
		end

reg Pass_688;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_688<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1833==mem[688])&&(Pass_687))
				Pass_688<=1;
			else
				Pass_688<=0;
		end

reg Pass_689;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_689<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1843==mem[689])&&(Pass_688))
				Pass_689<=1;
			else
				Pass_689<=0;
		end

reg Pass_690;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_690<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1853==mem[690])&&(Pass_689))
				Pass_690<=1;
			else
				Pass_690<=0;
		end

reg Pass_691;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_691<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1863==mem[691])&&(Pass_690))
				Pass_691<=1;
			else
				Pass_691<=0;
		end

reg Pass_692;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_692<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1873==mem[692])&&(Pass_691))
				Pass_692<=1;
			else
				Pass_692<=0;
		end

reg Pass_693;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_693<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1883==mem[693])&&(Pass_692))
				Pass_693<=1;
			else
				Pass_693<=0;
		end

reg Pass_694;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_694<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1893==mem[694])&&(Pass_693))
				Pass_694<=1;
			else
				Pass_694<=0;
		end

reg Pass_695;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_695<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18A3==mem[695])&&(Pass_694))
				Pass_695<=1;
			else
				Pass_695<=0;
		end

reg Pass_696;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_696<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18B3==mem[696])&&(Pass_695))
				Pass_696<=1;
			else
				Pass_696<=0;
		end

reg Pass_697;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_697<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18C3==mem[697])&&(Pass_696))
				Pass_697<=1;
			else
				Pass_697<=0;
		end

reg Pass_698;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_698<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18D3==mem[698])&&(Pass_697))
				Pass_698<=1;
			else
				Pass_698<=0;
		end

reg Pass_699;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_699<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P18E3==mem[699])&&(Pass_698))
				Pass_699<=1;
			else
				Pass_699<=0;
		end

reg Pass_700;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_700<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1913==mem[700])&&(Pass_699))
				Pass_700<=1;
			else
				Pass_700<=0;
		end

reg Pass_701;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_701<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1923==mem[701])&&(Pass_700))
				Pass_701<=1;
			else
				Pass_701<=0;
		end

reg Pass_702;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_702<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1933==mem[702])&&(Pass_701))
				Pass_702<=1;
			else
				Pass_702<=0;
		end

reg Pass_703;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_703<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1943==mem[703])&&(Pass_702))
				Pass_703<=1;
			else
				Pass_703<=0;
		end

reg Pass_704;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_704<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1953==mem[704])&&(Pass_703))
				Pass_704<=1;
			else
				Pass_704<=0;
		end

reg Pass_705;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_705<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1963==mem[705])&&(Pass_704))
				Pass_705<=1;
			else
				Pass_705<=0;
		end

reg Pass_706;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_706<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1973==mem[706])&&(Pass_705))
				Pass_706<=1;
			else
				Pass_706<=0;
		end

reg Pass_707;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_707<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1983==mem[707])&&(Pass_706))
				Pass_707<=1;
			else
				Pass_707<=0;
		end

reg Pass_708;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_708<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1993==mem[708])&&(Pass_707))
				Pass_708<=1;
			else
				Pass_708<=0;
		end

reg Pass_709;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_709<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19A3==mem[709])&&(Pass_708))
				Pass_709<=1;
			else
				Pass_709<=0;
		end

reg Pass_710;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_710<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19B3==mem[710])&&(Pass_709))
				Pass_710<=1;
			else
				Pass_710<=0;
		end

reg Pass_711;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_711<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19C3==mem[711])&&(Pass_710))
				Pass_711<=1;
			else
				Pass_711<=0;
		end

reg Pass_712;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_712<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19D3==mem[712])&&(Pass_711))
				Pass_712<=1;
			else
				Pass_712<=0;
		end

reg Pass_713;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_713<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P19E3==mem[713])&&(Pass_712))
				Pass_713<=1;
			else
				Pass_713<=0;
		end

reg Pass_714;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_714<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A13==mem[714])&&(Pass_713))
				Pass_714<=1;
			else
				Pass_714<=0;
		end

reg Pass_715;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_715<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A23==mem[715])&&(Pass_714))
				Pass_715<=1;
			else
				Pass_715<=0;
		end

reg Pass_716;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_716<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A33==mem[716])&&(Pass_715))
				Pass_716<=1;
			else
				Pass_716<=0;
		end

reg Pass_717;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_717<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A43==mem[717])&&(Pass_716))
				Pass_717<=1;
			else
				Pass_717<=0;
		end

reg Pass_718;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_718<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A53==mem[718])&&(Pass_717))
				Pass_718<=1;
			else
				Pass_718<=0;
		end

reg Pass_719;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_719<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A63==mem[719])&&(Pass_718))
				Pass_719<=1;
			else
				Pass_719<=0;
		end

reg Pass_720;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_720<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A73==mem[720])&&(Pass_719))
				Pass_720<=1;
			else
				Pass_720<=0;
		end

reg Pass_721;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_721<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A83==mem[721])&&(Pass_720))
				Pass_721<=1;
			else
				Pass_721<=0;
		end

reg Pass_722;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_722<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1A93==mem[722])&&(Pass_721))
				Pass_722<=1;
			else
				Pass_722<=0;
		end

reg Pass_723;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_723<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AA3==mem[723])&&(Pass_722))
				Pass_723<=1;
			else
				Pass_723<=0;
		end

reg Pass_724;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_724<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AB3==mem[724])&&(Pass_723))
				Pass_724<=1;
			else
				Pass_724<=0;
		end

reg Pass_725;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_725<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AC3==mem[725])&&(Pass_724))
				Pass_725<=1;
			else
				Pass_725<=0;
		end

reg Pass_726;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_726<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AD3==mem[726])&&(Pass_725))
				Pass_726<=1;
			else
				Pass_726<=0;
		end

reg Pass_727;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_727<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1AE3==mem[727])&&(Pass_726))
				Pass_727<=1;
			else
				Pass_727<=0;
		end

reg Pass_728;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_728<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B13==mem[728])&&(Pass_727))
				Pass_728<=1;
			else
				Pass_728<=0;
		end

reg Pass_729;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_729<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B23==mem[729])&&(Pass_728))
				Pass_729<=1;
			else
				Pass_729<=0;
		end

reg Pass_730;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_730<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B33==mem[730])&&(Pass_729))
				Pass_730<=1;
			else
				Pass_730<=0;
		end

reg Pass_731;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_731<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B43==mem[731])&&(Pass_730))
				Pass_731<=1;
			else
				Pass_731<=0;
		end

reg Pass_732;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_732<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B53==mem[732])&&(Pass_731))
				Pass_732<=1;
			else
				Pass_732<=0;
		end

reg Pass_733;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_733<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B63==mem[733])&&(Pass_732))
				Pass_733<=1;
			else
				Pass_733<=0;
		end

reg Pass_734;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_734<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B73==mem[734])&&(Pass_733))
				Pass_734<=1;
			else
				Pass_734<=0;
		end

reg Pass_735;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_735<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B83==mem[735])&&(Pass_734))
				Pass_735<=1;
			else
				Pass_735<=0;
		end

reg Pass_736;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_736<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1B93==mem[736])&&(Pass_735))
				Pass_736<=1;
			else
				Pass_736<=0;
		end

reg Pass_737;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_737<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BA3==mem[737])&&(Pass_736))
				Pass_737<=1;
			else
				Pass_737<=0;
		end

reg Pass_738;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_738<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BB3==mem[738])&&(Pass_737))
				Pass_738<=1;
			else
				Pass_738<=0;
		end

reg Pass_739;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_739<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BC3==mem[739])&&(Pass_738))
				Pass_739<=1;
			else
				Pass_739<=0;
		end

reg Pass_740;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_740<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BD3==mem[740])&&(Pass_739))
				Pass_740<=1;
			else
				Pass_740<=0;
		end

reg Pass_741;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_741<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1BE3==mem[741])&&(Pass_740))
				Pass_741<=1;
			else
				Pass_741<=0;
		end

reg Pass_742;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_742<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C13==mem[742])&&(Pass_741))
				Pass_742<=1;
			else
				Pass_742<=0;
		end

reg Pass_743;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_743<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C23==mem[743])&&(Pass_742))
				Pass_743<=1;
			else
				Pass_743<=0;
		end

reg Pass_744;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_744<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C33==mem[744])&&(Pass_743))
				Pass_744<=1;
			else
				Pass_744<=0;
		end

reg Pass_745;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_745<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C43==mem[745])&&(Pass_744))
				Pass_745<=1;
			else
				Pass_745<=0;
		end

reg Pass_746;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_746<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C53==mem[746])&&(Pass_745))
				Pass_746<=1;
			else
				Pass_746<=0;
		end

reg Pass_747;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_747<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C63==mem[747])&&(Pass_746))
				Pass_747<=1;
			else
				Pass_747<=0;
		end

reg Pass_748;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_748<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C73==mem[748])&&(Pass_747))
				Pass_748<=1;
			else
				Pass_748<=0;
		end

reg Pass_749;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_749<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C83==mem[749])&&(Pass_748))
				Pass_749<=1;
			else
				Pass_749<=0;
		end

reg Pass_750;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_750<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1C93==mem[750])&&(Pass_749))
				Pass_750<=1;
			else
				Pass_750<=0;
		end

reg Pass_751;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_751<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CA3==mem[751])&&(Pass_750))
				Pass_751<=1;
			else
				Pass_751<=0;
		end

reg Pass_752;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_752<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CB3==mem[752])&&(Pass_751))
				Pass_752<=1;
			else
				Pass_752<=0;
		end

reg Pass_753;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_753<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CC3==mem[753])&&(Pass_752))
				Pass_753<=1;
			else
				Pass_753<=0;
		end

reg Pass_754;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_754<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CD3==mem[754])&&(Pass_753))
				Pass_754<=1;
			else
				Pass_754<=0;
		end

reg Pass_755;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_755<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1CE3==mem[755])&&(Pass_754))
				Pass_755<=1;
			else
				Pass_755<=0;
		end

reg Pass_756;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_756<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D13==mem[756])&&(Pass_755))
				Pass_756<=1;
			else
				Pass_756<=0;
		end

reg Pass_757;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_757<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D23==mem[757])&&(Pass_756))
				Pass_757<=1;
			else
				Pass_757<=0;
		end

reg Pass_758;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_758<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D33==mem[758])&&(Pass_757))
				Pass_758<=1;
			else
				Pass_758<=0;
		end

reg Pass_759;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_759<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D43==mem[759])&&(Pass_758))
				Pass_759<=1;
			else
				Pass_759<=0;
		end

reg Pass_760;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_760<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D53==mem[760])&&(Pass_759))
				Pass_760<=1;
			else
				Pass_760<=0;
		end

reg Pass_761;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_761<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D63==mem[761])&&(Pass_760))
				Pass_761<=1;
			else
				Pass_761<=0;
		end

reg Pass_762;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_762<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D73==mem[762])&&(Pass_761))
				Pass_762<=1;
			else
				Pass_762<=0;
		end

reg Pass_763;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_763<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D83==mem[763])&&(Pass_762))
				Pass_763<=1;
			else
				Pass_763<=0;
		end

reg Pass_764;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_764<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1D93==mem[764])&&(Pass_763))
				Pass_764<=1;
			else
				Pass_764<=0;
		end

reg Pass_765;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_765<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DA3==mem[765])&&(Pass_764))
				Pass_765<=1;
			else
				Pass_765<=0;
		end

reg Pass_766;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_766<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DB3==mem[766])&&(Pass_765))
				Pass_766<=1;
			else
				Pass_766<=0;
		end

reg Pass_767;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_767<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DC3==mem[767])&&(Pass_766))
				Pass_767<=1;
			else
				Pass_767<=0;
		end

reg Pass_768;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_768<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DD3==mem[768])&&(Pass_767))
				Pass_768<=1;
			else
				Pass_768<=0;
		end

reg Pass_769;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_769<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1DE3==mem[769])&&(Pass_768))
				Pass_769<=1;
			else
				Pass_769<=0;
		end

reg Pass_770;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_770<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E13==mem[770])&&(Pass_769))
				Pass_770<=1;
			else
				Pass_770<=0;
		end

reg Pass_771;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_771<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E23==mem[771])&&(Pass_770))
				Pass_771<=1;
			else
				Pass_771<=0;
		end

reg Pass_772;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_772<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E33==mem[772])&&(Pass_771))
				Pass_772<=1;
			else
				Pass_772<=0;
		end

reg Pass_773;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_773<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E43==mem[773])&&(Pass_772))
				Pass_773<=1;
			else
				Pass_773<=0;
		end

reg Pass_774;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_774<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E53==mem[774])&&(Pass_773))
				Pass_774<=1;
			else
				Pass_774<=0;
		end

reg Pass_775;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_775<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E63==mem[775])&&(Pass_774))
				Pass_775<=1;
			else
				Pass_775<=0;
		end

reg Pass_776;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_776<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E73==mem[776])&&(Pass_775))
				Pass_776<=1;
			else
				Pass_776<=0;
		end

reg Pass_777;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_777<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E83==mem[777])&&(Pass_776))
				Pass_777<=1;
			else
				Pass_777<=0;
		end

reg Pass_778;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_778<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1E93==mem[778])&&(Pass_777))
				Pass_778<=1;
			else
				Pass_778<=0;
		end

reg Pass_779;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_779<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1EA3==mem[779])&&(Pass_778))
				Pass_779<=1;
			else
				Pass_779<=0;
		end

reg Pass_780;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_780<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1EB3==mem[780])&&(Pass_779))
				Pass_780<=1;
			else
				Pass_780<=0;
		end

reg Pass_781;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_781<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1EC3==mem[781])&&(Pass_780))
				Pass_781<=1;
			else
				Pass_781<=0;
		end

reg Pass_782;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_782<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1ED3==mem[782])&&(Pass_781))
				Pass_782<=1;
			else
				Pass_782<=0;
		end

reg Pass_783;
always@(posedge clk or negedge rstn)
	if(~rstn)
		Pass_783<=0;
	else if(count>=2)
		begin
			if((tb_test_layer0.test_layer0.P1EE3==mem[783])&&(Pass_782))
				Pass_783<=1;
			else
				Pass_783<=0;
		end

always@(posedge clk)
if(Pass_0&&Pass_1&&Pass_2&&Pass_3&&Pass_4&&Pass_5&&Pass_6&&Pass_7&&Pass_8&&Pass_9&&Pass_10&&Pass_11&&Pass_12&&Pass_13&&Pass_14&&Pass_15&&Pass_16&&Pass_17&&Pass_18&&Pass_19&&Pass_20&&Pass_21&&Pass_22&&Pass_23&&Pass_24&&Pass_25&&Pass_26&&Pass_27&&Pass_28&&Pass_29&&Pass_30&&Pass_31&&Pass_32&&Pass_33&&Pass_34&&Pass_35&&Pass_36&&Pass_37&&Pass_38&&Pass_39&&Pass_40&&Pass_41&&Pass_42&&Pass_43&&Pass_44&&Pass_45&&Pass_46&&Pass_47&&Pass_48&&Pass_49&&Pass_50&&Pass_51&&Pass_52&&Pass_53&&Pass_54&&Pass_55&&Pass_56&&Pass_57&&Pass_58&&Pass_59&&Pass_60&&Pass_61&&Pass_62&&Pass_63&&Pass_64&&Pass_65&&Pass_66&&Pass_67&&Pass_68&&Pass_69&&Pass_70&&Pass_71&&Pass_72&&Pass_73&&Pass_74&&Pass_75&&Pass_76&&Pass_77&&Pass_78&&Pass_79&&Pass_80&&Pass_81&&Pass_82&&Pass_83&&Pass_84&&Pass_85&&Pass_86&&Pass_87&&Pass_88&&Pass_89&&Pass_90&&Pass_91&&Pass_92&&Pass_93&&Pass_94&&Pass_95&&Pass_96&&Pass_97&&Pass_98&&Pass_99&&Pass_100&&Pass_101&&Pass_102&&Pass_103&&Pass_104&&Pass_105&&Pass_106&&Pass_107&&Pass_108&&Pass_109&&Pass_110&&Pass_111&&Pass_112&&Pass_113&&Pass_114&&Pass_115&&Pass_116&&Pass_117&&Pass_118&&Pass_119&&Pass_120&&Pass_121&&Pass_122&&Pass_123&&Pass_124&&Pass_125&&Pass_126&&Pass_127&&Pass_128&&Pass_129&&Pass_130&&Pass_131&&Pass_132&&Pass_133&&Pass_134&&Pass_135&&Pass_136&&Pass_137&&Pass_138&&Pass_139&&Pass_140&&Pass_141&&Pass_142&&Pass_143&&Pass_144&&Pass_145&&Pass_146&&Pass_147&&Pass_148&&Pass_149&&Pass_150&&Pass_151&&Pass_152&&Pass_153&&Pass_154&&Pass_155&&Pass_156&&Pass_157&&Pass_158&&Pass_159&&Pass_160&&Pass_161&&Pass_162&&Pass_163&&Pass_164&&Pass_165&&Pass_166&&Pass_167&&Pass_168&&Pass_169&&Pass_170&&Pass_171&&Pass_172&&Pass_173&&Pass_174&&Pass_175&&Pass_176&&Pass_177&&Pass_178&&Pass_179&&Pass_180&&Pass_181&&Pass_182&&Pass_183&&Pass_184&&Pass_185&&Pass_186&&Pass_187&&Pass_188&&Pass_189&&Pass_190&&Pass_191&&Pass_192&&Pass_193&&Pass_194&&Pass_195&&Pass_196&&Pass_197&&Pass_198&&Pass_199&&Pass_200&&Pass_201&&Pass_202&&Pass_203&&Pass_204&&Pass_205&&Pass_206&&Pass_207&&Pass_208&&Pass_209&&Pass_210&&Pass_211&&Pass_212&&Pass_213&&Pass_214&&Pass_215&&Pass_216&&Pass_217&&Pass_218&&Pass_219&&Pass_220&&Pass_221&&Pass_222&&Pass_223&&Pass_224&&Pass_225&&Pass_226&&Pass_227&&Pass_228&&Pass_229&&Pass_230&&Pass_231&&Pass_232&&Pass_233&&Pass_234&&Pass_235&&Pass_236&&Pass_237&&Pass_238&&Pass_239&&Pass_240&&Pass_241&&Pass_242&&Pass_243&&Pass_244&&Pass_245&&Pass_246&&Pass_247&&Pass_248&&Pass_249&&Pass_250&&Pass_251&&Pass_252&&Pass_253&&Pass_254&&Pass_255&&Pass_256&&Pass_257&&Pass_258&&Pass_259&&Pass_260&&Pass_261&&Pass_262&&Pass_263&&Pass_264&&Pass_265&&Pass_266&&Pass_267&&Pass_268&&Pass_269&&Pass_270&&Pass_271&&Pass_272&&Pass_273&&Pass_274&&Pass_275&&Pass_276&&Pass_277&&Pass_278&&Pass_279&&Pass_280&&Pass_281&&Pass_282&&Pass_283&&Pass_284&&Pass_285&&Pass_286&&Pass_287&&Pass_288&&Pass_289&&Pass_290&&Pass_291&&Pass_292&&Pass_293&&Pass_294&&Pass_295&&Pass_296&&Pass_297&&Pass_298&&Pass_299&&Pass_300&&Pass_301&&Pass_302&&Pass_303&&Pass_304&&Pass_305&&Pass_306&&Pass_307&&Pass_308&&Pass_309&&Pass_310&&Pass_311&&Pass_312&&Pass_313&&Pass_314&&Pass_315&&Pass_316&&Pass_317&&Pass_318&&Pass_319&&Pass_320&&Pass_321&&Pass_322&&Pass_323&&Pass_324&&Pass_325&&Pass_326&&Pass_327&&Pass_328&&Pass_329&&Pass_330&&Pass_331&&Pass_332&&Pass_333&&Pass_334&&Pass_335&&Pass_336&&Pass_337&&Pass_338&&Pass_339&&Pass_340&&Pass_341&&Pass_342&&Pass_343&&Pass_344&&Pass_345&&Pass_346&&Pass_347&&Pass_348&&Pass_349&&Pass_350&&Pass_351&&Pass_352&&Pass_353&&Pass_354&&Pass_355&&Pass_356&&Pass_357&&Pass_358&&Pass_359&&Pass_360&&Pass_361&&Pass_362&&Pass_363&&Pass_364&&Pass_365&&Pass_366&&Pass_367&&Pass_368&&Pass_369&&Pass_370&&Pass_371&&Pass_372&&Pass_373&&Pass_374&&Pass_375&&Pass_376&&Pass_377&&Pass_378&&Pass_379&&Pass_380&&Pass_381&&Pass_382&&Pass_383&&Pass_384&&Pass_385&&Pass_386&&Pass_387&&Pass_388&&Pass_389&&Pass_390&&Pass_391&&Pass_392&&Pass_393&&Pass_394&&Pass_395&&Pass_396&&Pass_397&&Pass_398&&Pass_399&&Pass_400&&Pass_401&&Pass_402&&Pass_403&&Pass_404&&Pass_405&&Pass_406&&Pass_407&&Pass_408&&Pass_409&&Pass_410&&Pass_411&&Pass_412&&Pass_413&&Pass_414&&Pass_415&&Pass_416&&Pass_417&&Pass_418&&Pass_419&&Pass_420&&Pass_421&&Pass_422&&Pass_423&&Pass_424&&Pass_425&&Pass_426&&Pass_427&&Pass_428&&Pass_429&&Pass_430&&Pass_431&&Pass_432&&Pass_433&&Pass_434&&Pass_435&&Pass_436&&Pass_437&&Pass_438&&Pass_439&&Pass_440&&Pass_441&&Pass_442&&Pass_443&&Pass_444&&Pass_445&&Pass_446&&Pass_447&&Pass_448&&Pass_449&&Pass_450&&Pass_451&&Pass_452&&Pass_453&&Pass_454&&Pass_455&&Pass_456&&Pass_457&&Pass_458&&Pass_459&&Pass_460&&Pass_461&&Pass_462&&Pass_463&&Pass_464&&Pass_465&&Pass_466&&Pass_467&&Pass_468&&Pass_469&&Pass_470&&Pass_471&&Pass_472&&Pass_473&&Pass_474&&Pass_475&&Pass_476&&Pass_477&&Pass_478&&Pass_479&&Pass_480&&Pass_481&&Pass_482&&Pass_483&&Pass_484&&Pass_485&&Pass_486&&Pass_487&&Pass_488&&Pass_489&&Pass_490&&Pass_491&&Pass_492&&Pass_493&&Pass_494&&Pass_495&&Pass_496&&Pass_497&&Pass_498&&Pass_499&&Pass_500&&Pass_501&&Pass_502&&Pass_503&&Pass_504&&Pass_505&&Pass_506&&Pass_507&&Pass_508&&Pass_509&&Pass_510&&Pass_511&&Pass_512&&Pass_513&&Pass_514&&Pass_515&&Pass_516&&Pass_517&&Pass_518&&Pass_519&&Pass_520&&Pass_521&&Pass_522&&Pass_523&&Pass_524&&Pass_525&&Pass_526&&Pass_527&&Pass_528&&Pass_529&&Pass_530&&Pass_531&&Pass_532&&Pass_533&&Pass_534&&Pass_535&&Pass_536&&Pass_537&&Pass_538&&Pass_539&&Pass_540&&Pass_541&&Pass_542&&Pass_543&&Pass_544&&Pass_545&&Pass_546&&Pass_547&&Pass_548&&Pass_549&&Pass_550&&Pass_551&&Pass_552&&Pass_553&&Pass_554&&Pass_555&&Pass_556&&Pass_557&&Pass_558&&Pass_559&&Pass_560&&Pass_561&&Pass_562&&Pass_563&&Pass_564&&Pass_565&&Pass_566&&Pass_567&&Pass_568&&Pass_569&&Pass_570&&Pass_571&&Pass_572&&Pass_573&&Pass_574&&Pass_575&&Pass_576&&Pass_577&&Pass_578&&Pass_579&&Pass_580&&Pass_581&&Pass_582&&Pass_583&&Pass_584&&Pass_585&&Pass_586&&Pass_587&&Pass_588&&Pass_589&&Pass_590&&Pass_591&&Pass_592&&Pass_593&&Pass_594&&Pass_595&&Pass_596&&Pass_597&&Pass_598&&Pass_599&&Pass_600&&Pass_601&&Pass_602&&Pass_603&&Pass_604&&Pass_605&&Pass_606&&Pass_607&&Pass_608&&Pass_609&&Pass_610&&Pass_611&&Pass_612&&Pass_613&&Pass_614&&Pass_615&&Pass_616&&Pass_617&&Pass_618&&Pass_619&&Pass_620&&Pass_621&&Pass_622&&Pass_623&&Pass_624&&Pass_625&&Pass_626&&Pass_627&&Pass_628&&Pass_629&&Pass_630&&Pass_631&&Pass_632&&Pass_633&&Pass_634&&Pass_635&&Pass_636&&Pass_637&&Pass_638&&Pass_639&&Pass_640&&Pass_641&&Pass_642&&Pass_643&&Pass_644&&Pass_645&&Pass_646&&Pass_647&&Pass_648&&Pass_649&&Pass_650&&Pass_651&&Pass_652&&Pass_653&&Pass_654&&Pass_655&&Pass_656&&Pass_657&&Pass_658&&Pass_659&&Pass_660&&Pass_661&&Pass_662&&Pass_663&&Pass_664&&Pass_665&&Pass_666&&Pass_667&&Pass_668&&Pass_669&&Pass_670&&Pass_671&&Pass_672&&Pass_673&&Pass_674&&Pass_675&&Pass_676&&Pass_677&&Pass_678&&Pass_679&&Pass_680&&Pass_681&&Pass_682&&Pass_683&&Pass_684&&Pass_685&&Pass_686&&Pass_687&&Pass_688&&Pass_689&&Pass_690&&Pass_691&&Pass_692&&Pass_693&&Pass_694&&Pass_695&&Pass_696&&Pass_697&&Pass_698&&Pass_699&&Pass_700&&Pass_701&&Pass_702&&Pass_703&&Pass_704&&Pass_705&&Pass_706&&Pass_707&&Pass_708&&Pass_709&&Pass_710&&Pass_711&&Pass_712&&Pass_713&&Pass_714&&Pass_715&&Pass_716&&Pass_717&&Pass_718&&Pass_719&&Pass_720&&Pass_721&&Pass_722&&Pass_723&&Pass_724&&Pass_725&&Pass_726&&Pass_727&&Pass_728&&Pass_729&&Pass_730&&Pass_731&&Pass_732&&Pass_733&&Pass_734&&Pass_735&&Pass_736&&Pass_737&&Pass_738&&Pass_739&&Pass_740&&Pass_741&&Pass_742&&Pass_743&&Pass_744&&Pass_745&&Pass_746&&Pass_747&&Pass_748&&Pass_749&&Pass_750&&Pass_751&&Pass_752&&Pass_753&&Pass_754&&Pass_755&&Pass_756&&Pass_757&&Pass_758&&Pass_759&&Pass_760&&Pass_761&&Pass_762&&Pass_763&&Pass_764&&Pass_765&&Pass_766&&Pass_767&&Pass_768&&Pass_769&&Pass_770&&Pass_771&&Pass_772&&Pass_773&&Pass_774&&Pass_775&&Pass_776&&Pass_777&&Pass_778&&Pass_779&&Pass_780&&Pass_781&&Pass_782&&Pass_783)
begin
$display("PASS");
$finish;
end

endmodule
